module AN2D0BWP16P90 (
	A1,
	A2,
	Z
);
	input wire A1;
	input wire A2;
	output wire Z;
	assign Z = A1 & A2;
endmodule
module AO22D0BWP16P90 (
	A1,
	A2,
	B1,
	B2,
	Z
);
	input wire A1;
	input wire A2;
	input wire B1;
	input wire B2;
	output wire Z;
	assign Z = (A1 & A2) | (B1 & B2);
endmodule
module sky130_sram_1kbyte_1rw1r_32x256_8 (
	clk0,
	csb0,
	web0,
	wmask0,
	addr0,
	din0,
	dout0,
	clk1,
	csb1,
	addr1,
	dout1
);
	parameter NUM_WMASKS = 4;
	parameter DATA_WIDTH = 32;
	parameter ADDR_WIDTH = 8;
	parameter RAM_DEPTH = 1 << ADDR_WIDTH;
	parameter DELAY = 0;
	input clk0;
	input csb0;
	input web0;
	input [NUM_WMASKS - 1:0] wmask0;
	input [ADDR_WIDTH - 1:0] addr0;
	input [DATA_WIDTH - 1:0] din0;
	output reg [DATA_WIDTH - 1:0] dout0;
	input clk1;
	input csb1;
	input [ADDR_WIDTH - 1:0] addr1;
	output reg [DATA_WIDTH - 1:0] dout1;
	reg csb0_reg;
	reg web0_reg;
	reg [NUM_WMASKS - 1:0] wmask0_reg;
	reg [ADDR_WIDTH - 1:0] addr0_reg;
	reg [DATA_WIDTH - 1:0] din0_reg;
	reg [DATA_WIDTH - 1:0] mem [0:RAM_DEPTH - 1];
	always @(posedge clk0) begin
		csb0_reg = csb0;
		web0_reg = web0;
		wmask0_reg = wmask0;
		addr0_reg = addr0;
		din0_reg = din0;
		//dout0 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	end
	reg csb1_reg;
	reg [ADDR_WIDTH - 1:0] addr1_reg;
	always @(posedge clk1) begin
		csb1_reg = csb1;
		addr1_reg = addr1;
		//dout1 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	end
	always @(negedge clk0) begin : MEM_WRITE0
		if (!csb0_reg && !web0_reg) begin
			if (wmask0_reg[0])
				mem[addr0_reg][7:0] = din0_reg[7:0];
			if (wmask0_reg[1])
				mem[addr0_reg][15:8] = din0_reg[15:8];
			if (wmask0_reg[2])
				mem[addr0_reg][23:16] = din0_reg[23:16];
			if (wmask0_reg[3])
				mem[addr0_reg][31:24] = din0_reg[31:24];
		end
	end
	always @(negedge clk0) begin : MEM_READ0
		if (!csb0_reg && web0_reg)
			dout0 <= #(DELAY) mem[addr0_reg];
	end
	always @(negedge clk1) begin : MEM_READ1
		if (!csb1_reg)
			dout1 <= #(DELAY) mem[addr1_reg];
	end
endmodule
module tile_en (
	I,
	O
);
	input [10:0] I;
	output [0:0] O;
	assign O = I[10];
endmodule
module mode (
	I,
	O
);
	input [10:0] I;
	output [1:0] O;
	assign O = I[9:8];
endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5 (
// 	I,
// 	O
// );
// 	input [10:0] I;
// 	output [3:0] O;
// 	assign O = I[7:4];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4 (
// 	I,
// 	O
// );
// 	input [10:0] I;
// 	output [3:0] O;
// 	assign O = I[3:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [3:0] O;
// 	assign O = I[31:28];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [3:0] O;
// 	assign O = I[27:24];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [3:0] O;
// 	assign O = I[23:20];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [3:0] O;
// 	assign O = I[19:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [3:0] O;
// 	assign O = I[15:12];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [3:0] O;
// 	assign O = I[11:8];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [3:0] O;
// 	assign O = I[7:4];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [3:0] O;
// 	assign O = I[3:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [3:0] O;
// 	assign O = I[31:28];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [3:0] O;
// 	assign O = I[27:24];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [3:0] O;
// 	assign O = I[23:20];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [3:0] O;
// 	assign O = I[19:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable (
// 	I,
// 	O
// );
// 	input [16:0] I;
// 	output [0:0] O;
// 	assign O = I[16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5 (
// 	I,
// 	O
// );
// 	input [16:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable (
// 	I,
// 	O
// );
// 	input [24:0] I;
// 	output [0:0] O;
// 	assign O = I[24];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5 (
// 	I,
// 	O
// );
// 	input [24:0] I;
// 	output [3:0] O;
// 	assign O = I[23:20];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4 (
// 	I,
// 	O
// );
// 	input [24:0] I;
// 	output [3:0] O;
// 	assign O = I[19:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3 (
// 	I,
// 	O
// );
// 	input [24:0] I;
// 	output [3:0] O;
// 	assign O = I[15:12];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2 (
// 	I,
// 	O
// );
// 	input [24:0] I;
// 	output [3:0] O;
// 	assign O = I[11:8];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1 (
// 	I,
// 	O
// );
// 	input [24:0] I;
// 	output [3:0] O;
// 	assign O = I[7:4];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0 (
// 	I,
// 	O
// );
// 	input [24:0] I;
// 	output [3:0] O;
// 	assign O = I[3:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [3:0] O;
// 	assign O = I[31:28];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [3:0] O;
// 	assign O = I[27:24];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [3:0] O;
// 	assign O = I[23:20];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [3:0] O;
// 	assign O = I[19:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [3:0] O;
// 	assign O = I[15:12];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [3:0] O;
// 	assign O = I[11:8];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [3:0] O;
// 	assign O = I[7:4];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [3:0] O;
// 	assign O = I[3:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality (
// 	I,
// 	O
// );
// 	input [19:0] I;
// 	output [3:0] O;
// 	assign O = I[19:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5 (
// 	I,
// 	O
// );
// 	input [19:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0 (
// 	I,
// 	O
// );
// 	input [19:0] I;
// 	output [15:0] O;
// 	assign O = I[19:4];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality (
// 	I,
// 	O
// );
// 	input [19:0] I;
// 	output [3:0] O;
// 	assign O = I[3:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr (
// 	I,
// 	O
// );
// 	input [16:0] I;
// 	output [15:0] O;
// 	assign O = I[16:1];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable (
// 	I,
// 	O
// );
// 	input [16:0] I;
// 	output [0:0] O;
// 	assign O = I[0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr (
// 	I,
// 	O
// );
// 	input [16:0] I;
// 	output [15:0] O;
// 	assign O = I[16:1];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable (
// 	I,
// 	O
// );
// 	input [16:0] I;
// 	output [0:0] O;
// 	assign O = I[0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality (
// 	I,
// 	O
// );
// 	input [19:0] I;
// 	output [3:0] O;
// 	assign O = I[19:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5 (
// 	I,
// 	O
// );
// 	input [19:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[31:16];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1 (
// 	I,
// 	O
// );
// 	input [31:0] I;
// 	output [15:0] O;
// 	assign O = I[15:0];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0 (
// 	I,
// 	O
// );
// 	input [27:0] I;
// 	output [15:0] O;
// 	assign O = I[27:12];
// endmodule
// module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality (
// 	I,
// 	O
// );
// 	input [27:0] I;
// 	output [3:0] O;
// 	assign O = I[11:8];
// endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5 (
	I,
	O
);
	input [27:0] I;
	output [7:0] O;
	assign O = I[7:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4 (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[31:24];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3 (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[23:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2 (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[15:8];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1 (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[7:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0 (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[31:24];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[23:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5 (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[15:8];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4 (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[7:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3 (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[31:24];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2 (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[23:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1 (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[15:8];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0 (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[7:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[31:24];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_5 (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[23:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_4 (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[15:8];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_3 (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[7:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_2 (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[31:24];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_1 (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[23:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_0 (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[15:8];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[7:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_5 (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[31:24];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_4 (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[23:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_3 (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[15:8];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_2 (
	I,
	O
);
	input [31:0] I;
	output [7:0] O;
	assign O = I[7:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_1 (
	I,
	O
);
	input [24:0] I;
	output [7:0] O;
	assign O = I[24:17];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_0 (
	I,
	O
);
	input [24:0] I;
	output [7:0] O;
	assign O = I[16:9];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr (
	I,
	O
);
	input [24:0] I;
	output [7:0] O;
	assign O = I[8:1];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en (
	I,
	O
);
	input [24:0] I;
	output [0:0] O;
	assign O = I[0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality (
	I,
	O
);
	input [19:0] I;
	output [3:0] O;
	assign O = I[19:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5 (
	I,
	O
);
	input [19:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0 (
	I,
	O
);
	input [19:0] I;
	output [15:0] O;
	assign O = I[19:4];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality (
	I,
	O
);
	input [19:0] I;
	output [3:0] O;
	assign O = I[3:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr (
	I,
	O
);
	input [16:0] I;
	output [15:0] O;
	assign O = I[16:1];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable (
	I,
	O
);
	input [16:0] I;
	output [0:0] O;
	assign O = I[0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr (
	I,
	O
);
	input [16:0] I;
	output [15:0] O;
	assign O = I[16:1];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable (
	I,
	O
);
	input [16:0] I;
	output [0:0] O;
	assign O = I[0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_5 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_4 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_3 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality (
	I,
	O
);
	input [19:0] I;
	output [3:0] O;
	assign O = I[19:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_5 (
	I,
	O
);
	input [19:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_4 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_3 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0 (
	I,
	O
);
	input [19:0] I;
	output [15:0] O;
	assign O = I[19:4];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality (
	I,
	O
);
	input [19:0] I;
	output [3:0] O;
	assign O = I[3:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr (
	I,
	O
);
	input [16:0] I;
	output [15:0] O;
	assign O = I[16:1];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable (
	I,
	O
);
	input [16:0] I;
	output [0:0] O;
	assign O = I[0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr (
	I,
	O
);
	input [16:0] I;
	output [15:0] O;
	assign O = I[16:1];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable (
	I,
	O
);
	input [16:0] I;
	output [0:0] O;
	assign O = I[0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_5 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[31:28];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_4 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[27:24];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_3 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[23:20];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[19:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[15:12];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[11:8];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[7:4];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_5 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[3:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_4 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[31:28];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_3 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[27:24];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[23:20];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[19:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[15:12];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[11:8];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_5 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[7:4];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_4 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[3:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_3 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[31:28];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_2 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[27:24];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_1 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[23:20];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_0 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[19:16];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[15:12];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_5 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[11:8];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_4 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[7:4];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_3 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[3:0];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_2 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[31:28];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_1 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[27:24];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_0 (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[23:20];
endmodule
module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr (
	I,
	O
);
	input [31:0] I;
	output [3:0] O;
	assign O = I[19:16];
endmodule
module mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable (
	I,
	O
);
	input [16:0] I;
	output [0:0] O;
	assign O = I[16];
endmodule
module mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5 (
	I,
	O
);
	input [16:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[31:16];
endmodule
module mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1 (
	I,
	O
);
	input [31:0] I;
	output [15:0] O;
	assign O = I[15:0];
endmodule
module mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0 (
	I,
	O
);
	input [25:0] I;
	output [15:0] O;
	assign O = I[25:10];
endmodule
module mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality (
	I,
	O
);
	input [25:0] I;
	output [3:0] O;
	assign O = I[9:6];
endmodule
module mantle_wire__typeBitIn9 (
	in,
	out
);
	output [8:0] in;
	input [8:0] out;
	assign in = out;
endmodule
module mantle_wire__typeBitIn8 (
	in,
	out
);
	output [7:0] in;
	input [7:0] out;
	assign in = out;
endmodule
module mantle_wire__typeBitIn7 (
	in,
	out
);
	output [6:0] in;
	input [6:0] out;
	assign in = out;
endmodule
module mantle_wire__typeBitIn67 (
	in,
	out
);
	output [66:0] in;
	input [66:0] out;
	assign in = out;
endmodule
module mantle_wire__typeBitIn4 (
	in,
	out
);
	output [3:0] in;
	input [3:0] out;
	assign in = out;
endmodule
module mantle_wire__typeBitIn32 (
	in,
	out
);
	output [31:0] in;
	input [31:0] out;
	assign in = out;
endmodule
module mantle_wire__typeBitIn3 (
	in,
	out
);
	output [2:0] in;
	input [2:0] out;
	assign in = out;
endmodule
module mantle_wire__typeBitIn2 (
	in,
	out
);
	output [1:0] in;
	input [1:0] out;
	assign in = out;
endmodule
module mantle_wire__typeBitIn16 (
	in,
	out
);
	output [15:0] in;
	input [15:0] out;
	assign in = out;
endmodule
module mantle_wire__typeBit9 (
	in,
	out
);
	input [8:0] in;
	output [8:0] out;
	assign out = in;
endmodule
module mantle_wire__typeBit8 (
	in,
	out
);
	input [7:0] in;
	output [7:0] out;
	assign out = in;
endmodule
module mantle_wire__typeBit4 (
	in,
	out
);
	input [3:0] in;
	output [3:0] out;
	assign out = in;
endmodule
module mantle_wire__typeBit32 (
	in,
	out
);
	input [31:0] in;
	output [31:0] out;
	assign out = in;
endmodule
module mantle_wire__typeBit30 (
	in,
	out
);
	input [29:0] in;
	output [29:0] out;
	assign out = in;
endmodule
module mantle_wire__typeBit28 (
	in,
	out
);
	input [27:0] in;
	output [27:0] out;
	assign out = in;
endmodule
module mantle_wire__typeBit26 (
	in,
	out
);
	input [25:0] in;
	output [25:0] out;
	assign out = in;
endmodule
module mantle_wire__typeBit25 (
	in,
	out
);
	input [24:0] in;
	output [24:0] out;
	assign out = in;
endmodule
module mantle_wire__typeBit20 (
	in,
	out
);
	input [19:0] in;
	output [19:0] out;
	assign out = in;
endmodule
module mantle_wire__typeBit18 (
	in,
	out
);
	input [17:0] in;
	output [17:0] out;
	assign out = in;
endmodule
module mantle_wire__typeBit17 (
	in,
	out
);
	input [16:0] in;
	output [16:0] out;
	assign out = in;
endmodule
module mantle_wire__typeBit16 (
	in,
	out
);
	input [15:0] in;
	output [15:0] out;
	assign out = in;
endmodule
module mantle_wire__typeBit11 (
	in,
	out
);
	input [10:0] in;
	output [10:0] out;
	assign out = in;
endmodule
module regCE_arst (
	in,
	ce,
	out,
	clk,
	arst
);
	parameter width = 1;
	parameter init = 1;
	input [width - 1:0] in;
	input ce;
	output [width - 1:0] out;
	input clk;
	input arst;
	reg [width - 1:0] value;
	always @(posedge clk or posedge arst)
		if (arst)
			value <= init;
		else if (ce)
			value <= in;
	assign out = value;
endmodule
module regCE (
	in,
	ce,
	out,
	clk
);
	parameter width = 1;
	input [width - 1:0] in;
	input ce;
	output [width - 1:0] out;
	input clk;
	reg [width - 1:0] value;
	always @(posedge clk)
		if (ce)
			value <= in;
	assign out = value;
endmodule
module io_core (
	glb2io_16,
	glb2io_1,
	io2glb_16,
	io2glb_1,
	f2io_16,
	f2io_1,
	io2f_16,
	io2f_1
);
	input [15:0] glb2io_16;
	input [0:0] glb2io_1;
	output [15:0] io2glb_16;
	output [0:0] io2glb_1;
	input [15:0] f2io_16;
	input [0:0] f2io_1;
	output [15:0] io2f_16;
	output [0:0] io2f_1;
	assign io2glb_16 = f2io_16;
	assign io2glb_1 = f2io_1;
	assign io2f_16 = glb2io_16;
	assign io2f_1 = glb2io_1;
endmodule
module inst_2 (
	I,
	O
);
	input [31:0] I;
	output [31:0] O;
	assign O = I;
endmodule
module inst_1 (
	I,
	O
);
	input [31:0] I;
	output [31:0] O;
	assign O = I;
endmodule
module inst_0 (
	I,
	O
);
	input [31:0] I;
	output [31:0] O;
	assign O = I;
endmodule
module input_width_1_num_1_reg_value (
	I,
	O
);
	input [25:0] I;
	output [0:0] O;
	assign O = I[5];
endmodule
module input_width_1_num_1_reg_sel (
	I,
	O
);
	input [25:0] I;
	output [0:0] O;
	assign O = I[4];
endmodule
module input_width_1_num_0_reg_value (
	I,
	O
);
	input [25:0] I;
	output [0:0] O;
	assign O = I[3];
endmodule
module input_width_1_num_0_reg_sel (
	I,
	O
);
	input [25:0] I;
	output [0:0] O;
	assign O = I[2];
endmodule
module flush_reg_value (
	I,
	O
);
	input [25:0] I;
	output [0:0] O;
	assign O = I[1];
endmodule
module flush_reg_sel (
	I,
	O
);
	input [25:0] I;
	output [0:0] O;
	assign O = I[0];
endmodule
module coreir_xor (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output [width - 1:0] out;
	assign out = in0 ^ in1;
endmodule
module coreir_wrap (
	in,
	out
);
	input in;
	output out;
	assign out = in;
endmodule
module coreir_ult (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output out;
	assign out = in0 < in1;
endmodule
module coreir_ule (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output out;
	assign out = in0 <= in1;
endmodule
module coreir_ugt (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output out;
	assign out = in0 > in1;
endmodule
module coreir_uge (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output out;
	assign out = in0 >= in1;
endmodule
module coreir_sub (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output [width - 1:0] out;
	assign out = in0 - in1;
endmodule
module coreir_slt (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output out;
	assign out = $signed(in0) < $signed(in1);
endmodule
module coreir_slice (
	in,
	out
);
	parameter hi = 1;
	parameter lo = 0;
	parameter width = 1;
	input [width - 1:0] in;
	output [(hi - lo) - 1:0] out;
	assign out = in[hi - 1:lo];
endmodule
module coreir_sle (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output out;
	assign out = $signed(in0) <= $signed(in1);
endmodule
module coreir_shl (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output [width - 1:0] out;
	assign out = in0 << in1;
endmodule
module coreir_sge (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output out;
	assign out = $signed(in0) >= $signed(in1);
endmodule
module coreir_reg_arst (
	clk,
	arst,
	in,
	out
);
	parameter width = 1;
	parameter arst_posedge = 1;
	parameter clk_posedge = 1;
	parameter init = 1;
	input clk;
	input arst;
	input [width - 1:0] in;
	output [width - 1:0] out;
	reg [width - 1:0] outReg;
	wire real_rst;
	assign real_rst = (arst_posedge ? arst : ~arst);
	wire real_clk;
	assign real_clk = (clk_posedge ? clk : ~clk);
	always @(posedge real_clk or posedge real_rst)
		if (real_rst)
			outReg <= init;
		else
			outReg <= in;
	assign out = outReg;
endmodule
module coreir_orr (
	in,
	out
);
	parameter width = 1;
	input [width - 1:0] in;
	output out;
	assign out = |in;
endmodule
module coreir_or (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output [width - 1:0] out;
	assign out = in0 | in1;
endmodule
module coreir_not (
	in,
	out
);
	parameter width = 1;
	input [width - 1:0] in;
	output [width - 1:0] out;
	assign out = ~in;
endmodule
module coreir_neg (
	in,
	out
);
	parameter width = 1;
	input [width - 1:0] in;
	output [width - 1:0] out;
	assign out = -in;
endmodule
module coreir_mux (
	in0,
	in1,
	sel,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	input sel;
	output [width - 1:0] out;
	assign out = (sel ? in1 : in0);
endmodule
module coreir_mul (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output [width - 1:0] out;
	assign out = in0 * in1;
endmodule
module coreir_lshr (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output [width - 1:0] out;
	assign out = in0 >> in1;
endmodule
module coreir_eq (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output out;
	assign out = in0 == in1;
endmodule
module coreir_const (out);
	parameter width = 1;
	parameter value = 1;
	output [width - 1:0] out;
	assign out = value;
endmodule
module coreir_ashr (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output [width - 1:0] out;
	assign out = $signed(in0) >>> in1;
endmodule
module coreir_and (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output [width - 1:0] out;
	assign out = in0 & in1;
endmodule
module coreir_add (
	in0,
	in1,
	out
);
	parameter width = 1;
	input [width - 1:0] in0;
	input [width - 1:0] in1;
	output [width - 1:0] out;
	assign out = in0 + in1;
endmodule
module corebit_xor (
	in0,
	in1,
	out
);
	input in0;
	input in1;
	output out;
	assign out = in0 ^ in1;
endmodule
module corebit_term (in);
	input in;
endmodule
module corebit_or (
	in0,
	in1,
	out
);
	input in0;
	input in1;
	output out;
	assign out = in0 | in1;
endmodule
module corebit_not (
	in,
	out
);
	input in;
	output out;
	assign out = ~in;
endmodule
module corebit_const (out);
	parameter value = 1;
	output out;
	assign out = value;
endmodule
module corebit_and (
	in0,
	in1,
	out
);
	input in0;
	input in1;
	output out;
	assign out = in0 & in1;
endmodule
module commonlib_muxn__N2__width32 (
	in_data_0,
	in_data_1,
	in_sel,
	out
);
	input [31:0] in_data_0;
	input [31:0] in_data_1;
	input [0:0] in_sel;
	output [31:0] out;
	wire [31:0] _join_out;
	coreir_mux #(.width(32)) _join(
		.in0(in_data_0),
		.in1(in_data_1),
		.sel(in_sel[0]),
		.out(_join_out)
	);
	assign out = _join_out;
endmodule
module commonlib_muxn__N4__width32 (
	in_data_0,
	in_data_1,
	in_data_2,
	in_data_3,
	in_sel,
	out
);
	input [31:0] in_data_0;
	input [31:0] in_data_1;
	input [31:0] in_data_2;
	input [31:0] in_data_3;
	input [1:0] in_sel;
	output [31:0] out;
	wire [31:0] _join_out;
	wire [31:0] muxN_0_out;
	wire [31:0] muxN_1_out;
	wire [0:0] sel_slice0_out;
	wire [0:0] sel_slice1_out;
	coreir_mux #(.width(32)) _join(
		.in0(muxN_0_out),
		.in1(muxN_1_out),
		.sel(in_sel[1]),
		.out(_join_out)
	);
	commonlib_muxn__N2__width32 muxN_0(
		.in_data_0(in_data_0),
		.in_data_1(in_data_1),
		.in_sel(sel_slice0_out),
		.out(muxN_0_out)
	);
	commonlib_muxn__N2__width32 muxN_1(
		.in_data_0(in_data_2),
		.in_data_1(in_data_3),
		.in_sel(sel_slice1_out),
		.out(muxN_1_out)
	);
	coreir_slice #(
		.hi(1),
		.lo(0),
		.width(2)
	) sel_slice0(
		.in(in_sel),
		.out(sel_slice0_out)
	);
	coreir_slice #(
		.hi(1),
		.lo(0),
		.width(2)
	) sel_slice1(
		.in(in_sel),
		.out(sel_slice1_out)
	);
	assign out = _join_out;
endmodule
module commonlib_muxn__N8__width32 (
	in_data_0,
	in_data_1,
	in_data_2,
	in_data_3,
	in_data_4,
	in_data_5,
	in_data_6,
	in_data_7,
	in_sel,
	out
);
	input [31:0] in_data_0;
	input [31:0] in_data_1;
	input [31:0] in_data_2;
	input [31:0] in_data_3;
	input [31:0] in_data_4;
	input [31:0] in_data_5;
	input [31:0] in_data_6;
	input [31:0] in_data_7;
	input [2:0] in_sel;
	output [31:0] out;
	wire [31:0] _join_out;
	wire [31:0] muxN_0_out;
	wire [31:0] muxN_1_out;
	wire [1:0] sel_slice0_out;
	wire [1:0] sel_slice1_out;
	coreir_mux #(.width(32)) _join(
		.in0(muxN_0_out),
		.in1(muxN_1_out),
		.sel(in_sel[2]),
		.out(_join_out)
	);
	commonlib_muxn__N4__width32 muxN_0(
		.in_data_0(in_data_0),
		.in_data_1(in_data_1),
		.in_data_2(in_data_2),
		.in_data_3(in_data_3),
		.in_sel(sel_slice0_out),
		.out(muxN_0_out)
	);
	commonlib_muxn__N4__width32 muxN_1(
		.in_data_0(in_data_4),
		.in_data_1(in_data_5),
		.in_data_2(in_data_6),
		.in_data_3(in_data_7),
		.in_sel(sel_slice1_out),
		.out(muxN_1_out)
	);
	coreir_slice #(
		.hi(2),
		.lo(0),
		.width(3)
	) sel_slice0(
		.in(in_sel),
		.out(sel_slice0_out)
	);
	coreir_slice #(
		.hi(2),
		.lo(0),
		.width(3)
	) sel_slice1(
		.in(in_sel),
		.out(sel_slice1_out)
	);
	assign out = _join_out;
endmodule
module commonlib_muxn__N2__width16 (
	in_data_0,
	in_data_1,
	in_sel,
	out
);
	input [15:0] in_data_0;
	input [15:0] in_data_1;
	input [0:0] in_sel;
	output [15:0] out;
	wire [15:0] _join_out;
	coreir_mux #(.width(16)) _join(
		.in0(in_data_0),
		.in1(in_data_1),
		.sel(in_sel[0]),
		.out(_join_out)
	);
	assign out = _join_out;
endmodule
module commonlib_muxn__N4__width16 (
	in_data_0,
	in_data_1,
	in_data_2,
	in_data_3,
	in_sel,
	out
);
	input [15:0] in_data_0;
	input [15:0] in_data_1;
	input [15:0] in_data_2;
	input [15:0] in_data_3;
	input [1:0] in_sel;
	output [15:0] out;
	wire [15:0] _join_out;
	wire [15:0] muxN_0_out;
	wire [15:0] muxN_1_out;
	wire [0:0] sel_slice0_out;
	wire [0:0] sel_slice1_out;
	coreir_mux #(.width(16)) _join(
		.in0(muxN_0_out),
		.in1(muxN_1_out),
		.sel(in_sel[1]),
		.out(_join_out)
	);
	commonlib_muxn__N2__width16 muxN_0(
		.in_data_0(in_data_0),
		.in_data_1(in_data_1),
		.in_sel(sel_slice0_out),
		.out(muxN_0_out)
	);
	commonlib_muxn__N2__width16 muxN_1(
		.in_data_0(in_data_2),
		.in_data_1(in_data_3),
		.in_sel(sel_slice1_out),
		.out(muxN_1_out)
	);
	coreir_slice #(
		.hi(1),
		.lo(0),
		.width(2)
	) sel_slice0(
		.in(in_sel),
		.out(sel_slice0_out)
	);
	coreir_slice #(
		.hi(1),
		.lo(0),
		.width(2)
	) sel_slice1(
		.in(in_sel),
		.out(sel_slice1_out)
	);
	assign out = _join_out;
endmodule
module commonlib_muxn__N8__width16 (
	in_data_0,
	in_data_1,
	in_data_2,
	in_data_3,
	in_data_4,
	in_data_5,
	in_data_6,
	in_data_7,
	in_sel,
	out
);
	input [15:0] in_data_0;
	input [15:0] in_data_1;
	input [15:0] in_data_2;
	input [15:0] in_data_3;
	input [15:0] in_data_4;
	input [15:0] in_data_5;
	input [15:0] in_data_6;
	input [15:0] in_data_7;
	input [2:0] in_sel;
	output [15:0] out;
	wire [15:0] _join_out;
	wire [15:0] muxN_0_out;
	wire [15:0] muxN_1_out;
	wire [1:0] sel_slice0_out;
	wire [1:0] sel_slice1_out;
	coreir_mux #(.width(16)) _join(
		.in0(muxN_0_out),
		.in1(muxN_1_out),
		.sel(in_sel[2]),
		.out(_join_out)
	);
	commonlib_muxn__N4__width16 muxN_0(
		.in_data_0(in_data_0),
		.in_data_1(in_data_1),
		.in_data_2(in_data_2),
		.in_data_3(in_data_3),
		.in_sel(sel_slice0_out),
		.out(muxN_0_out)
	);
	commonlib_muxn__N4__width16 muxN_1(
		.in_data_0(in_data_4),
		.in_data_1(in_data_5),
		.in_data_2(in_data_6),
		.in_data_3(in_data_7),
		.in_sel(sel_slice1_out),
		.out(muxN_1_out)
	);
	coreir_slice #(
		.hi(2),
		.lo(0),
		.width(3)
	) sel_slice0(
		.in(in_sel),
		.out(sel_slice0_out)
	);
	coreir_slice #(
		.hi(2),
		.lo(0),
		.width(3)
	) sel_slice1(
		.in(in_sel),
		.out(sel_slice1_out)
	);
	assign out = _join_out;
endmodule
module commonlib_muxn__N2__width1 (
	in_data_0,
	in_data_1,
	in_sel,
	out
);
	input [0:0] in_data_0;
	input [0:0] in_data_1;
	input [0:0] in_sel;
	output [0:0] out;
	wire [0:0] _join_out;
	coreir_mux #(.width(1)) _join(
		.in0(in_data_0),
		.in1(in_data_1),
		.sel(in_sel[0]),
		.out(_join_out)
	);
	assign out = _join_out;
endmodule
module commonlib_muxn__N4__width1 (
	in_data_0,
	in_data_1,
	in_data_2,
	in_data_3,
	in_sel,
	out
);
	input [0:0] in_data_0;
	input [0:0] in_data_1;
	input [0:0] in_data_2;
	input [0:0] in_data_3;
	input [1:0] in_sel;
	output [0:0] out;
	wire [0:0] _join_out;
	wire [0:0] muxN_0_out;
	wire [0:0] muxN_1_out;
	wire [0:0] sel_slice0_out;
	wire [0:0] sel_slice1_out;
	coreir_mux #(.width(1)) _join(
		.in0(muxN_0_out),
		.in1(muxN_1_out),
		.sel(in_sel[1]),
		.out(_join_out)
	);
	commonlib_muxn__N2__width1 muxN_0(
		.in_data_0(in_data_0),
		.in_data_1(in_data_1),
		.in_sel(sel_slice0_out),
		.out(muxN_0_out)
	);
	commonlib_muxn__N2__width1 muxN_1(
		.in_data_0(in_data_2),
		.in_data_1(in_data_3),
		.in_sel(sel_slice1_out),
		.out(muxN_1_out)
	);
	coreir_slice #(
		.hi(1),
		.lo(0),
		.width(2)
	) sel_slice0(
		.in(in_sel),
		.out(sel_slice0_out)
	);
	coreir_slice #(
		.hi(1),
		.lo(0),
		.width(2)
	) sel_slice1(
		.in(in_sel),
		.out(sel_slice1_out)
	);
	assign out = _join_out;
endmodule
module commonlib_muxn__N8__width1 (
	in_data_0,
	in_data_1,
	in_data_2,
	in_data_3,
	in_data_4,
	in_data_5,
	in_data_6,
	in_data_7,
	in_sel,
	out
);
	input [0:0] in_data_0;
	input [0:0] in_data_1;
	input [0:0] in_data_2;
	input [0:0] in_data_3;
	input [0:0] in_data_4;
	input [0:0] in_data_5;
	input [0:0] in_data_6;
	input [0:0] in_data_7;
	input [2:0] in_sel;
	output [0:0] out;
	wire [0:0] _join_out;
	wire [0:0] muxN_0_out;
	wire [0:0] muxN_1_out;
	wire [1:0] sel_slice0_out;
	wire [1:0] sel_slice1_out;
	coreir_mux #(.width(1)) _join(
		.in0(muxN_0_out),
		.in1(muxN_1_out),
		.sel(in_sel[2]),
		.out(_join_out)
	);
	commonlib_muxn__N4__width1 muxN_0(
		.in_data_0(in_data_0),
		.in_data_1(in_data_1),
		.in_data_2(in_data_2),
		.in_data_3(in_data_3),
		.in_sel(sel_slice0_out),
		.out(muxN_0_out)
	);
	commonlib_muxn__N4__width1 muxN_1(
		.in_data_0(in_data_4),
		.in_data_1(in_data_5),
		.in_data_2(in_data_6),
		.in_data_3(in_data_7),
		.in_sel(sel_slice1_out),
		.out(muxN_1_out)
	);
	coreir_slice #(
		.hi(2),
		.lo(0),
		.width(3)
	) sel_slice0(
		.in(in_sel),
		.out(sel_slice0_out)
	);
	coreir_slice #(
		.hi(2),
		.lo(0),
		.width(3)
	) sel_slice1(
		.in(in_sel),
		.out(sel_slice1_out)
	);
	assign out = _join_out;
endmodule
module commonlib_muxn__N6__width1 (
	in_data_0,
	in_data_1,
	in_data_2,
	in_data_3,
	in_data_4,
	in_data_5,
	in_sel,
	out
);
	input [0:0] in_data_0;
	input [0:0] in_data_1;
	input [0:0] in_data_2;
	input [0:0] in_data_3;
	input [0:0] in_data_4;
	input [0:0] in_data_5;
	input [2:0] in_sel;
	output [0:0] out;
	wire [0:0] _join_out;
	wire [0:0] muxN_0_out;
	wire [0:0] muxN_1_out;
	wire [1:0] sel_slice0_out;
	wire [0:0] sel_slice1_out;
	coreir_mux #(.width(1)) _join(
		.in0(muxN_0_out),
		.in1(muxN_1_out),
		.sel(in_sel[2]),
		.out(_join_out)
	);
	commonlib_muxn__N4__width1 muxN_0(
		.in_data_0(in_data_0),
		.in_data_1(in_data_1),
		.in_data_2(in_data_2),
		.in_data_3(in_data_3),
		.in_sel(sel_slice0_out),
		.out(muxN_0_out)
	);
	commonlib_muxn__N2__width1 muxN_1(
		.in_data_0(in_data_4),
		.in_data_1(in_data_5),
		.in_sel(sel_slice1_out),
		.out(muxN_1_out)
	);
	coreir_slice #(
		.hi(2),
		.lo(0),
		.width(3)
	) sel_slice0(
		.in(in_sel),
		.out(sel_slice0_out)
	);
	coreir_slice #(
		.hi(1),
		.lo(0),
		.width(3)
	) sel_slice1(
		.in(in_sel),
		.out(sel_slice1_out)
	);
	assign out = _join_out;
endmodule
module commonlib_muxn__N1__width32 (
	in_data_0,
	in_sel,
	out
);
	input [31:0] in_data_0;
	input [0:0] in_sel;
	output [31:0] out;
	corebit_term term_sel(.in(in_sel[0]));
	assign out = in_data_0;
endmodule
module commonlib_muxn__N3__width32 (
	in_data_0,
	in_data_1,
	in_data_2,
	in_sel,
	out
);
	input [31:0] in_data_0;
	input [31:0] in_data_1;
	input [31:0] in_data_2;
	input [1:0] in_sel;
	output [31:0] out;
	wire [31:0] _join_out;
	wire [31:0] muxN_0_out;
	wire [31:0] muxN_1_out;
	wire [0:0] sel_slice0_out;
	wire [0:0] sel_slice1_out;
	coreir_mux #(.width(32)) _join(
		.in0(muxN_0_out),
		.in1(muxN_1_out),
		.sel(in_sel[1]),
		.out(_join_out)
	);
	commonlib_muxn__N2__width32 muxN_0(
		.in_data_0(in_data_0),
		.in_data_1(in_data_1),
		.in_sel(sel_slice0_out),
		.out(muxN_0_out)
	);
	commonlib_muxn__N1__width32 muxN_1(
		.in_data_0(in_data_2),
		.in_sel(sel_slice1_out),
		.out(muxN_1_out)
	);
	coreir_slice #(
		.hi(1),
		.lo(0),
		.width(2)
	) sel_slice0(
		.in(in_sel),
		.out(sel_slice0_out)
	);
	coreir_slice #(
		.hi(1),
		.lo(0),
		.width(2)
	) sel_slice1(
		.in(in_sel),
		.out(sel_slice1_out)
	);
	assign out = _join_out;
endmodule
module commonlib_muxn__N1__width16 (
	in_data_0,
	in_sel,
	out
);
	input [15:0] in_data_0;
	input [0:0] in_sel;
	output [15:0] out;
	corebit_term term_sel(.in(in_sel[0]));
	assign out = in_data_0;
endmodule
module commonlib_muxn__N5__width16 (
	in_data_0,
	in_data_1,
	in_data_2,
	in_data_3,
	in_data_4,
	in_sel,
	out
);
	input [15:0] in_data_0;
	input [15:0] in_data_1;
	input [15:0] in_data_2;
	input [15:0] in_data_3;
	input [15:0] in_data_4;
	input [2:0] in_sel;
	output [15:0] out;
	wire [15:0] _join_out;
	wire [15:0] muxN_0_out;
	wire [15:0] muxN_1_out;
	wire [1:0] sel_slice0_out;
	wire [0:0] sel_slice1_out;
	coreir_mux #(.width(16)) _join(
		.in0(muxN_0_out),
		.in1(muxN_1_out),
		.sel(in_sel[2]),
		.out(_join_out)
	);
	commonlib_muxn__N4__width16 muxN_0(
		.in_data_0(in_data_0),
		.in_data_1(in_data_1),
		.in_data_2(in_data_2),
		.in_data_3(in_data_3),
		.in_sel(sel_slice0_out),
		.out(muxN_0_out)
	);
	commonlib_muxn__N1__width16 muxN_1(
		.in_data_0(in_data_4),
		.in_sel(sel_slice1_out),
		.out(muxN_1_out)
	);
	coreir_slice #(
		.hi(2),
		.lo(0),
		.width(3)
	) sel_slice0(
		.in(in_sel),
		.out(sel_slice0_out)
	);
	coreir_slice #(
		.hi(1),
		.lo(0),
		.width(3)
	) sel_slice1(
		.in(in_sel),
		.out(sel_slice1_out)
	);
	assign out = _join_out;
endmodule
module commonlib_muxn__N16__width32 (
	in_data_0,
	in_data_1,
	in_data_10,
	in_data_11,
	in_data_12,
	in_data_13,
	in_data_14,
	in_data_15,
	in_data_2,
	in_data_3,
	in_data_4,
	in_data_5,
	in_data_6,
	in_data_7,
	in_data_8,
	in_data_9,
	in_sel,
	out
);
	input [31:0] in_data_0;
	input [31:0] in_data_1;
	input [31:0] in_data_10;
	input [31:0] in_data_11;
	input [31:0] in_data_12;
	input [31:0] in_data_13;
	input [31:0] in_data_14;
	input [31:0] in_data_15;
	input [31:0] in_data_2;
	input [31:0] in_data_3;
	input [31:0] in_data_4;
	input [31:0] in_data_5;
	input [31:0] in_data_6;
	input [31:0] in_data_7;
	input [31:0] in_data_8;
	input [31:0] in_data_9;
	input [3:0] in_sel;
	output [31:0] out;
	wire [31:0] _join_out;
	wire [31:0] muxN_0_out;
	wire [31:0] muxN_1_out;
	wire [2:0] sel_slice0_out;
	wire [2:0] sel_slice1_out;
	coreir_mux #(.width(32)) _join(
		.in0(muxN_0_out),
		.in1(muxN_1_out),
		.sel(in_sel[3]),
		.out(_join_out)
	);
	commonlib_muxn__N8__width32 muxN_0(
		.in_data_0(in_data_0),
		.in_data_1(in_data_1),
		.in_data_2(in_data_2),
		.in_data_3(in_data_3),
		.in_data_4(in_data_4),
		.in_data_5(in_data_5),
		.in_data_6(in_data_6),
		.in_data_7(in_data_7),
		.in_sel(sel_slice0_out),
		.out(muxN_0_out)
	);
	commonlib_muxn__N8__width32 muxN_1(
		.in_data_0(in_data_8),
		.in_data_1(in_data_9),
		.in_data_2(in_data_10),
		.in_data_3(in_data_11),
		.in_data_4(in_data_12),
		.in_data_5(in_data_13),
		.in_data_6(in_data_14),
		.in_data_7(in_data_15),
		.in_sel(sel_slice1_out),
		.out(muxN_1_out)
	);
	coreir_slice #(
		.hi(3),
		.lo(0),
		.width(4)
	) sel_slice0(
		.in(in_sel),
		.out(sel_slice0_out)
	);
	coreir_slice #(
		.hi(3),
		.lo(0),
		.width(4)
	) sel_slice1(
		.in(in_sel),
		.out(sel_slice1_out)
	);
	assign out = _join_out;
endmodule
module commonlib_muxn__N32__width32 (
	in_data_0,
	in_data_1,
	in_data_10,
	in_data_11,
	in_data_12,
	in_data_13,
	in_data_14,
	in_data_15,
	in_data_16,
	in_data_17,
	in_data_18,
	in_data_19,
	in_data_2,
	in_data_20,
	in_data_21,
	in_data_22,
	in_data_23,
	in_data_24,
	in_data_25,
	in_data_26,
	in_data_27,
	in_data_28,
	in_data_29,
	in_data_3,
	in_data_30,
	in_data_31,
	in_data_4,
	in_data_5,
	in_data_6,
	in_data_7,
	in_data_8,
	in_data_9,
	in_sel,
	out
);
	input [31:0] in_data_0;
	input [31:0] in_data_1;
	input [31:0] in_data_10;
	input [31:0] in_data_11;
	input [31:0] in_data_12;
	input [31:0] in_data_13;
	input [31:0] in_data_14;
	input [31:0] in_data_15;
	input [31:0] in_data_16;
	input [31:0] in_data_17;
	input [31:0] in_data_18;
	input [31:0] in_data_19;
	input [31:0] in_data_2;
	input [31:0] in_data_20;
	input [31:0] in_data_21;
	input [31:0] in_data_22;
	input [31:0] in_data_23;
	input [31:0] in_data_24;
	input [31:0] in_data_25;
	input [31:0] in_data_26;
	input [31:0] in_data_27;
	input [31:0] in_data_28;
	input [31:0] in_data_29;
	input [31:0] in_data_3;
	input [31:0] in_data_30;
	input [31:0] in_data_31;
	input [31:0] in_data_4;
	input [31:0] in_data_5;
	input [31:0] in_data_6;
	input [31:0] in_data_7;
	input [31:0] in_data_8;
	input [31:0] in_data_9;
	input [4:0] in_sel;
	output [31:0] out;
	wire [31:0] _join_out;
	wire [31:0] muxN_0_out;
	wire [31:0] muxN_1_out;
	wire [3:0] sel_slice0_out;
	wire [3:0] sel_slice1_out;
	coreir_mux #(.width(32)) _join(
		.in0(muxN_0_out),
		.in1(muxN_1_out),
		.sel(in_sel[4]),
		.out(_join_out)
	);
	commonlib_muxn__N16__width32 muxN_0(
		.in_data_0(in_data_0),
		.in_data_1(in_data_1),
		.in_data_10(in_data_10),
		.in_data_11(in_data_11),
		.in_data_12(in_data_12),
		.in_data_13(in_data_13),
		.in_data_14(in_data_14),
		.in_data_15(in_data_15),
		.in_data_2(in_data_2),
		.in_data_3(in_data_3),
		.in_data_4(in_data_4),
		.in_data_5(in_data_5),
		.in_data_6(in_data_6),
		.in_data_7(in_data_7),
		.in_data_8(in_data_8),
		.in_data_9(in_data_9),
		.in_sel(sel_slice0_out),
		.out(muxN_0_out)
	);
	commonlib_muxn__N16__width32 muxN_1(
		.in_data_0(in_data_16),
		.in_data_1(in_data_17),
		.in_data_10(in_data_26),
		.in_data_11(in_data_27),
		.in_data_12(in_data_28),
		.in_data_13(in_data_29),
		.in_data_14(in_data_30),
		.in_data_15(in_data_31),
		.in_data_2(in_data_18),
		.in_data_3(in_data_19),
		.in_data_4(in_data_20),
		.in_data_5(in_data_21),
		.in_data_6(in_data_22),
		.in_data_7(in_data_23),
		.in_data_8(in_data_24),
		.in_data_9(in_data_25),
		.in_sel(sel_slice1_out),
		.out(muxN_1_out)
	);
	coreir_slice #(
		.hi(4),
		.lo(0),
		.width(5)
	) sel_slice0(
		.in(in_sel),
		.out(sel_slice0_out)
	);
	coreir_slice #(
		.hi(4),
		.lo(0),
		.width(5)
	) sel_slice1(
		.in(in_sel),
		.out(sel_slice1_out)
	);
	assign out = _join_out;
endmodule
module commonlib_muxn__N64__width32 (
	in_data_0,
	in_data_1,
	in_data_10,
	in_data_11,
	in_data_12,
	in_data_13,
	in_data_14,
	in_data_15,
	in_data_16,
	in_data_17,
	in_data_18,
	in_data_19,
	in_data_2,
	in_data_20,
	in_data_21,
	in_data_22,
	in_data_23,
	in_data_24,
	in_data_25,
	in_data_26,
	in_data_27,
	in_data_28,
	in_data_29,
	in_data_3,
	in_data_30,
	in_data_31,
	in_data_32,
	in_data_33,
	in_data_34,
	in_data_35,
	in_data_36,
	in_data_37,
	in_data_38,
	in_data_39,
	in_data_4,
	in_data_40,
	in_data_41,
	in_data_42,
	in_data_43,
	in_data_44,
	in_data_45,
	in_data_46,
	in_data_47,
	in_data_48,
	in_data_49,
	in_data_5,
	in_data_50,
	in_data_51,
	in_data_52,
	in_data_53,
	in_data_54,
	in_data_55,
	in_data_56,
	in_data_57,
	in_data_58,
	in_data_59,
	in_data_6,
	in_data_60,
	in_data_61,
	in_data_62,
	in_data_63,
	in_data_7,
	in_data_8,
	in_data_9,
	in_sel,
	out
);
	input [31:0] in_data_0;
	input [31:0] in_data_1;
	input [31:0] in_data_10;
	input [31:0] in_data_11;
	input [31:0] in_data_12;
	input [31:0] in_data_13;
	input [31:0] in_data_14;
	input [31:0] in_data_15;
	input [31:0] in_data_16;
	input [31:0] in_data_17;
	input [31:0] in_data_18;
	input [31:0] in_data_19;
	input [31:0] in_data_2;
	input [31:0] in_data_20;
	input [31:0] in_data_21;
	input [31:0] in_data_22;
	input [31:0] in_data_23;
	input [31:0] in_data_24;
	input [31:0] in_data_25;
	input [31:0] in_data_26;
	input [31:0] in_data_27;
	input [31:0] in_data_28;
	input [31:0] in_data_29;
	input [31:0] in_data_3;
	input [31:0] in_data_30;
	input [31:0] in_data_31;
	input [31:0] in_data_32;
	input [31:0] in_data_33;
	input [31:0] in_data_34;
	input [31:0] in_data_35;
	input [31:0] in_data_36;
	input [31:0] in_data_37;
	input [31:0] in_data_38;
	input [31:0] in_data_39;
	input [31:0] in_data_4;
	input [31:0] in_data_40;
	input [31:0] in_data_41;
	input [31:0] in_data_42;
	input [31:0] in_data_43;
	input [31:0] in_data_44;
	input [31:0] in_data_45;
	input [31:0] in_data_46;
	input [31:0] in_data_47;
	input [31:0] in_data_48;
	input [31:0] in_data_49;
	input [31:0] in_data_5;
	input [31:0] in_data_50;
	input [31:0] in_data_51;
	input [31:0] in_data_52;
	input [31:0] in_data_53;
	input [31:0] in_data_54;
	input [31:0] in_data_55;
	input [31:0] in_data_56;
	input [31:0] in_data_57;
	input [31:0] in_data_58;
	input [31:0] in_data_59;
	input [31:0] in_data_6;
	input [31:0] in_data_60;
	input [31:0] in_data_61;
	input [31:0] in_data_62;
	input [31:0] in_data_63;
	input [31:0] in_data_7;
	input [31:0] in_data_8;
	input [31:0] in_data_9;
	input [5:0] in_sel;
	output [31:0] out;
	wire [31:0] _join_out;
	wire [31:0] muxN_0_out;
	wire [31:0] muxN_1_out;
	wire [4:0] sel_slice0_out;
	wire [4:0] sel_slice1_out;
	coreir_mux #(.width(32)) _join(
		.in0(muxN_0_out),
		.in1(muxN_1_out),
		.sel(in_sel[5]),
		.out(_join_out)
	);
	commonlib_muxn__N32__width32 muxN_0(
		.in_data_0(in_data_0),
		.in_data_1(in_data_1),
		.in_data_10(in_data_10),
		.in_data_11(in_data_11),
		.in_data_12(in_data_12),
		.in_data_13(in_data_13),
		.in_data_14(in_data_14),
		.in_data_15(in_data_15),
		.in_data_16(in_data_16),
		.in_data_17(in_data_17),
		.in_data_18(in_data_18),
		.in_data_19(in_data_19),
		.in_data_2(in_data_2),
		.in_data_20(in_data_20),
		.in_data_21(in_data_21),
		.in_data_22(in_data_22),
		.in_data_23(in_data_23),
		.in_data_24(in_data_24),
		.in_data_25(in_data_25),
		.in_data_26(in_data_26),
		.in_data_27(in_data_27),
		.in_data_28(in_data_28),
		.in_data_29(in_data_29),
		.in_data_3(in_data_3),
		.in_data_30(in_data_30),
		.in_data_31(in_data_31),
		.in_data_4(in_data_4),
		.in_data_5(in_data_5),
		.in_data_6(in_data_6),
		.in_data_7(in_data_7),
		.in_data_8(in_data_8),
		.in_data_9(in_data_9),
		.in_sel(sel_slice0_out),
		.out(muxN_0_out)
	);
	commonlib_muxn__N32__width32 muxN_1(
		.in_data_0(in_data_32),
		.in_data_1(in_data_33),
		.in_data_10(in_data_42),
		.in_data_11(in_data_43),
		.in_data_12(in_data_44),
		.in_data_13(in_data_45),
		.in_data_14(in_data_46),
		.in_data_15(in_data_47),
		.in_data_16(in_data_48),
		.in_data_17(in_data_49),
		.in_data_18(in_data_50),
		.in_data_19(in_data_51),
		.in_data_2(in_data_34),
		.in_data_20(in_data_52),
		.in_data_21(in_data_53),
		.in_data_22(in_data_54),
		.in_data_23(in_data_55),
		.in_data_24(in_data_56),
		.in_data_25(in_data_57),
		.in_data_26(in_data_58),
		.in_data_27(in_data_59),
		.in_data_28(in_data_60),
		.in_data_29(in_data_61),
		.in_data_3(in_data_35),
		.in_data_30(in_data_62),
		.in_data_31(in_data_63),
		.in_data_4(in_data_36),
		.in_data_5(in_data_37),
		.in_data_6(in_data_38),
		.in_data_7(in_data_39),
		.in_data_8(in_data_40),
		.in_data_9(in_data_41),
		.in_sel(sel_slice1_out),
		.out(muxN_1_out)
	);
	coreir_slice #(
		.hi(5),
		.lo(0),
		.width(6)
	) sel_slice0(
		.in(in_sel),
		.out(sel_slice0_out)
	);
	coreir_slice #(
		.hi(5),
		.lo(0),
		.width(6)
	) sel_slice1(
		.in(in_sel),
		.out(sel_slice1_out)
	);
	assign out = _join_out;
endmodule
module commonlib_muxn__N18__width32 (
	in_data_0,
	in_data_1,
	in_data_10,
	in_data_11,
	in_data_12,
	in_data_13,
	in_data_14,
	in_data_15,
	in_data_16,
	in_data_17,
	in_data_2,
	in_data_3,
	in_data_4,
	in_data_5,
	in_data_6,
	in_data_7,
	in_data_8,
	in_data_9,
	in_sel,
	out
);
	input [31:0] in_data_0;
	input [31:0] in_data_1;
	input [31:0] in_data_10;
	input [31:0] in_data_11;
	input [31:0] in_data_12;
	input [31:0] in_data_13;
	input [31:0] in_data_14;
	input [31:0] in_data_15;
	input [31:0] in_data_16;
	input [31:0] in_data_17;
	input [31:0] in_data_2;
	input [31:0] in_data_3;
	input [31:0] in_data_4;
	input [31:0] in_data_5;
	input [31:0] in_data_6;
	input [31:0] in_data_7;
	input [31:0] in_data_8;
	input [31:0] in_data_9;
	input [4:0] in_sel;
	output [31:0] out;
	wire [31:0] _join_out;
	wire [31:0] muxN_0_out;
	wire [31:0] muxN_1_out;
	wire [3:0] sel_slice0_out;
	wire [0:0] sel_slice1_out;
	coreir_mux #(.width(32)) _join(
		.in0(muxN_0_out),
		.in1(muxN_1_out),
		.sel(in_sel[4]),
		.out(_join_out)
	);
	commonlib_muxn__N16__width32 muxN_0(
		.in_data_0(in_data_0),
		.in_data_1(in_data_1),
		.in_data_10(in_data_10),
		.in_data_11(in_data_11),
		.in_data_12(in_data_12),
		.in_data_13(in_data_13),
		.in_data_14(in_data_14),
		.in_data_15(in_data_15),
		.in_data_2(in_data_2),
		.in_data_3(in_data_3),
		.in_data_4(in_data_4),
		.in_data_5(in_data_5),
		.in_data_6(in_data_6),
		.in_data_7(in_data_7),
		.in_data_8(in_data_8),
		.in_data_9(in_data_9),
		.in_sel(sel_slice0_out),
		.out(muxN_0_out)
	);
	commonlib_muxn__N2__width32 muxN_1(
		.in_data_0(in_data_16),
		.in_data_1(in_data_17),
		.in_sel(sel_slice1_out),
		.out(muxN_1_out)
	);
	coreir_slice #(
		.hi(4),
		.lo(0),
		.width(5)
	) sel_slice0(
		.in(in_sel),
		.out(sel_slice0_out)
	);
	coreir_slice #(
		.hi(1),
		.lo(0),
		.width(5)
	) sel_slice1(
		.in(in_sel),
		.out(sel_slice1_out)
	);
	assign out = _join_out;
endmodule
module commonlib_muxn__N82__width32 (
	in_data_0,
	in_data_1,
	in_data_10,
	in_data_11,
	in_data_12,
	in_data_13,
	in_data_14,
	in_data_15,
	in_data_16,
	in_data_17,
	in_data_18,
	in_data_19,
	in_data_2,
	in_data_20,
	in_data_21,
	in_data_22,
	in_data_23,
	in_data_24,
	in_data_25,
	in_data_26,
	in_data_27,
	in_data_28,
	in_data_29,
	in_data_3,
	in_data_30,
	in_data_31,
	in_data_32,
	in_data_33,
	in_data_34,
	in_data_35,
	in_data_36,
	in_data_37,
	in_data_38,
	in_data_39,
	in_data_4,
	in_data_40,
	in_data_41,
	in_data_42,
	in_data_43,
	in_data_44,
	in_data_45,
	in_data_46,
	in_data_47,
	in_data_48,
	in_data_49,
	in_data_5,
	in_data_50,
	in_data_51,
	in_data_52,
	in_data_53,
	in_data_54,
	in_data_55,
	in_data_56,
	in_data_57,
	in_data_58,
	in_data_59,
	in_data_6,
	in_data_60,
	in_data_61,
	in_data_62,
	in_data_63,
	in_data_64,
	in_data_65,
	in_data_66,
	in_data_67,
	in_data_68,
	in_data_69,
	in_data_7,
	in_data_70,
	in_data_71,
	in_data_72,
	in_data_73,
	in_data_74,
	in_data_75,
	in_data_76,
	in_data_77,
	in_data_78,
	in_data_79,
	in_data_8,
	in_data_80,
	in_data_81,
	in_data_9,
	in_sel,
	out
);
	input [31:0] in_data_0;
	input [31:0] in_data_1;
	input [31:0] in_data_10;
	input [31:0] in_data_11;
	input [31:0] in_data_12;
	input [31:0] in_data_13;
	input [31:0] in_data_14;
	input [31:0] in_data_15;
	input [31:0] in_data_16;
	input [31:0] in_data_17;
	input [31:0] in_data_18;
	input [31:0] in_data_19;
	input [31:0] in_data_2;
	input [31:0] in_data_20;
	input [31:0] in_data_21;
	input [31:0] in_data_22;
	input [31:0] in_data_23;
	input [31:0] in_data_24;
	input [31:0] in_data_25;
	input [31:0] in_data_26;
	input [31:0] in_data_27;
	input [31:0] in_data_28;
	input [31:0] in_data_29;
	input [31:0] in_data_3;
	input [31:0] in_data_30;
	input [31:0] in_data_31;
	input [31:0] in_data_32;
	input [31:0] in_data_33;
	input [31:0] in_data_34;
	input [31:0] in_data_35;
	input [31:0] in_data_36;
	input [31:0] in_data_37;
	input [31:0] in_data_38;
	input [31:0] in_data_39;
	input [31:0] in_data_4;
	input [31:0] in_data_40;
	input [31:0] in_data_41;
	input [31:0] in_data_42;
	input [31:0] in_data_43;
	input [31:0] in_data_44;
	input [31:0] in_data_45;
	input [31:0] in_data_46;
	input [31:0] in_data_47;
	input [31:0] in_data_48;
	input [31:0] in_data_49;
	input [31:0] in_data_5;
	input [31:0] in_data_50;
	input [31:0] in_data_51;
	input [31:0] in_data_52;
	input [31:0] in_data_53;
	input [31:0] in_data_54;
	input [31:0] in_data_55;
	input [31:0] in_data_56;
	input [31:0] in_data_57;
	input [31:0] in_data_58;
	input [31:0] in_data_59;
	input [31:0] in_data_6;
	input [31:0] in_data_60;
	input [31:0] in_data_61;
	input [31:0] in_data_62;
	input [31:0] in_data_63;
	input [31:0] in_data_64;
	input [31:0] in_data_65;
	input [31:0] in_data_66;
	input [31:0] in_data_67;
	input [31:0] in_data_68;
	input [31:0] in_data_69;
	input [31:0] in_data_7;
	input [31:0] in_data_70;
	input [31:0] in_data_71;
	input [31:0] in_data_72;
	input [31:0] in_data_73;
	input [31:0] in_data_74;
	input [31:0] in_data_75;
	input [31:0] in_data_76;
	input [31:0] in_data_77;
	input [31:0] in_data_78;
	input [31:0] in_data_79;
	input [31:0] in_data_8;
	input [31:0] in_data_80;
	input [31:0] in_data_81;
	input [31:0] in_data_9;
	input [6:0] in_sel;
	output [31:0] out;
	wire [31:0] _join_out;
	wire [31:0] muxN_0_out;
	wire [31:0] muxN_1_out;
	wire [5:0] sel_slice0_out;
	wire [4:0] sel_slice1_out;
	coreir_mux #(.width(32)) _join(
		.in0(muxN_0_out),
		.in1(muxN_1_out),
		.sel(in_sel[6]),
		.out(_join_out)
	);
	commonlib_muxn__N64__width32 muxN_0(
		.in_data_0(in_data_0),
		.in_data_1(in_data_1),
		.in_data_10(in_data_10),
		.in_data_11(in_data_11),
		.in_data_12(in_data_12),
		.in_data_13(in_data_13),
		.in_data_14(in_data_14),
		.in_data_15(in_data_15),
		.in_data_16(in_data_16),
		.in_data_17(in_data_17),
		.in_data_18(in_data_18),
		.in_data_19(in_data_19),
		.in_data_2(in_data_2),
		.in_data_20(in_data_20),
		.in_data_21(in_data_21),
		.in_data_22(in_data_22),
		.in_data_23(in_data_23),
		.in_data_24(in_data_24),
		.in_data_25(in_data_25),
		.in_data_26(in_data_26),
		.in_data_27(in_data_27),
		.in_data_28(in_data_28),
		.in_data_29(in_data_29),
		.in_data_3(in_data_3),
		.in_data_30(in_data_30),
		.in_data_31(in_data_31),
		.in_data_32(in_data_32),
		.in_data_33(in_data_33),
		.in_data_34(in_data_34),
		.in_data_35(in_data_35),
		.in_data_36(in_data_36),
		.in_data_37(in_data_37),
		.in_data_38(in_data_38),
		.in_data_39(in_data_39),
		.in_data_4(in_data_4),
		.in_data_40(in_data_40),
		.in_data_41(in_data_41),
		.in_data_42(in_data_42),
		.in_data_43(in_data_43),
		.in_data_44(in_data_44),
		.in_data_45(in_data_45),
		.in_data_46(in_data_46),
		.in_data_47(in_data_47),
		.in_data_48(in_data_48),
		.in_data_49(in_data_49),
		.in_data_5(in_data_5),
		.in_data_50(in_data_50),
		.in_data_51(in_data_51),
		.in_data_52(in_data_52),
		.in_data_53(in_data_53),
		.in_data_54(in_data_54),
		.in_data_55(in_data_55),
		.in_data_56(in_data_56),
		.in_data_57(in_data_57),
		.in_data_58(in_data_58),
		.in_data_59(in_data_59),
		.in_data_6(in_data_6),
		.in_data_60(in_data_60),
		.in_data_61(in_data_61),
		.in_data_62(in_data_62),
		.in_data_63(in_data_63),
		.in_data_7(in_data_7),
		.in_data_8(in_data_8),
		.in_data_9(in_data_9),
		.in_sel(sel_slice0_out),
		.out(muxN_0_out)
	);
	commonlib_muxn__N18__width32 muxN_1(
		.in_data_0(in_data_64),
		.in_data_1(in_data_65),
		.in_data_10(in_data_74),
		.in_data_11(in_data_75),
		.in_data_12(in_data_76),
		.in_data_13(in_data_77),
		.in_data_14(in_data_78),
		.in_data_15(in_data_79),
		.in_data_16(in_data_80),
		.in_data_17(in_data_81),
		.in_data_2(in_data_66),
		.in_data_3(in_data_67),
		.in_data_4(in_data_68),
		.in_data_5(in_data_69),
		.in_data_6(in_data_70),
		.in_data_7(in_data_71),
		.in_data_8(in_data_72),
		.in_data_9(in_data_73),
		.in_sel(sel_slice1_out),
		.out(muxN_1_out)
	);
	coreir_slice #(
		.hi(6),
		.lo(0),
		.width(7)
	) sel_slice0(
		.in(in_sel),
		.out(sel_slice0_out)
	);
	coreir_slice #(
		.hi(5),
		.lo(0),
		.width(7)
	) sel_slice1(
		.in(in_sel),
		.out(sel_slice1_out)
	);
	assign out = _join_out;
endmodule
module commonlib_muxn__N12__width16 (
	in_data_0,
	in_data_1,
	in_data_10,
	in_data_11,
	in_data_2,
	in_data_3,
	in_data_4,
	in_data_5,
	in_data_6,
	in_data_7,
	in_data_8,
	in_data_9,
	in_sel,
	out
);
	input [15:0] in_data_0;
	input [15:0] in_data_1;
	input [15:0] in_data_10;
	input [15:0] in_data_11;
	input [15:0] in_data_2;
	input [15:0] in_data_3;
	input [15:0] in_data_4;
	input [15:0] in_data_5;
	input [15:0] in_data_6;
	input [15:0] in_data_7;
	input [15:0] in_data_8;
	input [15:0] in_data_9;
	input [3:0] in_sel;
	output [15:0] out;
	wire [15:0] _join_out;
	wire [15:0] muxN_0_out;
	wire [15:0] muxN_1_out;
	wire [2:0] sel_slice0_out;
	wire [1:0] sel_slice1_out;
	coreir_mux #(.width(16)) _join(
		.in0(muxN_0_out),
		.in1(muxN_1_out),
		.sel(in_sel[3]),
		.out(_join_out)
	);
	commonlib_muxn__N8__width16 muxN_0(
		.in_data_0(in_data_0),
		.in_data_1(in_data_1),
		.in_data_2(in_data_2),
		.in_data_3(in_data_3),
		.in_data_4(in_data_4),
		.in_data_5(in_data_5),
		.in_data_6(in_data_6),
		.in_data_7(in_data_7),
		.in_sel(sel_slice0_out),
		.out(muxN_0_out)
	);
	commonlib_muxn__N4__width16 muxN_1(
		.in_data_0(in_data_8),
		.in_data_1(in_data_9),
		.in_data_2(in_data_10),
		.in_data_3(in_data_11),
		.in_sel(sel_slice1_out),
		.out(muxN_1_out)
	);
	coreir_slice #(
		.hi(3),
		.lo(0),
		.width(4)
	) sel_slice0(
		.in(in_sel),
		.out(sel_slice0_out)
	);
	coreir_slice #(
		.hi(2),
		.lo(0),
		.width(4)
	) sel_slice1(
		.in(in_sel),
		.out(sel_slice1_out)
	);
	assign out = _join_out;
endmodule
module commonlib_muxn__N12__width1 (
	in_data_0,
	in_data_1,
	in_data_10,
	in_data_11,
	in_data_2,
	in_data_3,
	in_data_4,
	in_data_5,
	in_data_6,
	in_data_7,
	in_data_8,
	in_data_9,
	in_sel,
	out
);
	input [0:0] in_data_0;
	input [0:0] in_data_1;
	input [0:0] in_data_10;
	input [0:0] in_data_11;
	input [0:0] in_data_2;
	input [0:0] in_data_3;
	input [0:0] in_data_4;
	input [0:0] in_data_5;
	input [0:0] in_data_6;
	input [0:0] in_data_7;
	input [0:0] in_data_8;
	input [0:0] in_data_9;
	input [3:0] in_sel;
	output [0:0] out;
	wire [0:0] _join_out;
	wire [0:0] muxN_0_out;
	wire [0:0] muxN_1_out;
	wire [2:0] sel_slice0_out;
	wire [1:0] sel_slice1_out;
	coreir_mux #(.width(1)) _join(
		.in0(muxN_0_out),
		.in1(muxN_1_out),
		.sel(in_sel[3]),
		.out(_join_out)
	);
	commonlib_muxn__N8__width1 muxN_0(
		.in_data_0(in_data_0),
		.in_data_1(in_data_1),
		.in_data_2(in_data_2),
		.in_data_3(in_data_3),
		.in_data_4(in_data_4),
		.in_data_5(in_data_5),
		.in_data_6(in_data_6),
		.in_data_7(in_data_7),
		.in_sel(sel_slice0_out),
		.out(muxN_0_out)
	);
	commonlib_muxn__N4__width1 muxN_1(
		.in_data_0(in_data_8),
		.in_data_1(in_data_9),
		.in_data_2(in_data_10),
		.in_data_3(in_data_11),
		.in_sel(sel_slice1_out),
		.out(muxN_1_out)
	);
	coreir_slice #(
		.hi(3),
		.lo(0),
		.width(4)
	) sel_slice0(
		.in(in_sel),
		.out(sel_slice0_out)
	);
	coreir_slice #(
		.hi(2),
		.lo(0),
		.width(4)
	) sel_slice1(
		.in(in_sel),
		.out(sel_slice1_out)
	);
	assign out = _join_out;
endmodule
module commonlib_muxn__N11__width32 (
	in_data_0,
	in_data_1,
	in_data_10,
	in_data_2,
	in_data_3,
	in_data_4,
	in_data_5,
	in_data_6,
	in_data_7,
	in_data_8,
	in_data_9,
	in_sel,
	out
);
	input [31:0] in_data_0;
	input [31:0] in_data_1;
	input [31:0] in_data_10;
	input [31:0] in_data_2;
	input [31:0] in_data_3;
	input [31:0] in_data_4;
	input [31:0] in_data_5;
	input [31:0] in_data_6;
	input [31:0] in_data_7;
	input [31:0] in_data_8;
	input [31:0] in_data_9;
	input [3:0] in_sel;
	output [31:0] out;
	wire [31:0] _join_out;
	wire [31:0] muxN_0_out;
	wire [31:0] muxN_1_out;
	wire [2:0] sel_slice0_out;
	wire [1:0] sel_slice1_out;
	coreir_mux #(.width(32)) _join(
		.in0(muxN_0_out),
		.in1(muxN_1_out),
		.sel(in_sel[3]),
		.out(_join_out)
	);
	commonlib_muxn__N8__width32 muxN_0(
		.in_data_0(in_data_0),
		.in_data_1(in_data_1),
		.in_data_2(in_data_2),
		.in_data_3(in_data_3),
		.in_data_4(in_data_4),
		.in_data_5(in_data_5),
		.in_data_6(in_data_6),
		.in_data_7(in_data_7),
		.in_sel(sel_slice0_out),
		.out(muxN_0_out)
	);
	commonlib_muxn__N3__width32 muxN_1(
		.in_data_0(in_data_8),
		.in_data_1(in_data_9),
		.in_data_2(in_data_10),
		.in_sel(sel_slice1_out),
		.out(muxN_1_out)
	);
	coreir_slice #(
		.hi(3),
		.lo(0),
		.width(4)
	) sel_slice0(
		.in(in_sel),
		.out(sel_slice0_out)
	);
	coreir_slice #(
		.hi(2),
		.lo(0),
		.width(4)
	) sel_slice1(
		.in(in_sel),
		.out(sel_slice1_out)
	);
	assign out = _join_out;
endmodule
module SB_T2_WEST_SB_OUT_B1_sel_unq1 (
	I,
	O
);
	input [17:0] I;
	output [2:0] O;
	assign O = I[17:15];
endmodule
module SB_T2_WEST_SB_OUT_B1_sel (
	I,
	O
);
	input [3:0] I;
	output [1:0] O;
	assign O = I[3:2];
endmodule
module SB_T2_WEST_SB_OUT_B16_sel_unq1 (
	I,
	O
);
	input [17:0] I;
	output [2:0] O;
	assign O = I[17:15];
endmodule
module SB_T2_WEST_SB_OUT_B16_sel (
	I,
	O
);
	input [3:0] I;
	output [1:0] O;
	assign O = I[3:2];
endmodule
module SB_T2_SOUTH_SB_OUT_B1_sel_unq1 (
	I,
	O
);
	input [17:0] I;
	output [2:0] O;
	assign O = I[14:12];
endmodule
module SB_T2_SOUTH_SB_OUT_B1_sel (
	I,
	O
);
	input [3:0] I;
	output [1:0] O;
	assign O = I[1:0];
endmodule
module SB_T2_SOUTH_SB_OUT_B16_sel_unq1 (
	I,
	O
);
	input [17:0] I;
	output [2:0] O;
	assign O = I[14:12];
endmodule
module SB_T2_SOUTH_SB_OUT_B16_sel (
	I,
	O
);
	input [3:0] I;
	output [1:0] O;
	assign O = I[1:0];
endmodule
module SB_T2_NORTH_SB_OUT_B1_sel_unq1 (
	I,
	O
);
	input [17:0] I;
	output [2:0] O;
	assign O = I[11:9];
endmodule
module SB_T2_NORTH_SB_OUT_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [1:0] O;
	assign O = I[31:30];
endmodule
module SB_T2_NORTH_SB_OUT_B16_sel_unq1 (
	I,
	O
);
	input [17:0] I;
	output [2:0] O;
	assign O = I[11:9];
endmodule
module SB_T2_NORTH_SB_OUT_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [1:0] O;
	assign O = I[31:30];
endmodule
module SB_T2_EAST_SB_OUT_B1_sel_unq1 (
	I,
	O
);
	input [17:0] I;
	output [2:0] O;
	assign O = I[8:6];
endmodule
module SB_T2_EAST_SB_OUT_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [1:0] O;
	assign O = I[29:28];
endmodule
module SB_T2_EAST_SB_OUT_B16_sel_unq1 (
	I,
	O
);
	input [17:0] I;
	output [2:0] O;
	assign O = I[8:6];
endmodule
module SB_T2_EAST_SB_OUT_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [1:0] O;
	assign O = I[29:28];
endmodule
module SB_T1_WEST_SB_OUT_B1_sel_unq1 (
	I,
	O
);
	input [17:0] I;
	output [2:0] O;
	assign O = I[5:3];
endmodule
module SB_T1_WEST_SB_OUT_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [1:0] O;
	assign O = I[27:26];
endmodule
module SB_T1_WEST_SB_OUT_B16_sel_unq1 (
	I,
	O
);
	input [17:0] I;
	output [2:0] O;
	assign O = I[5:3];
endmodule
module SB_T1_WEST_SB_OUT_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [1:0] O;
	assign O = I[27:26];
endmodule
module SB_T1_SOUTH_SB_OUT_B1_sel_unq1 (
	I,
	O
);
	input [17:0] I;
	output [2:0] O;
	assign O = I[2:0];
endmodule
module SB_T1_SOUTH_SB_OUT_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [1:0] O;
	assign O = I[25:24];
endmodule
module SB_T1_SOUTH_SB_OUT_B16_sel_unq1 (
	I,
	O
);
	input [17:0] I;
	output [2:0] O;
	assign O = I[2:0];
endmodule
module SB_T1_SOUTH_SB_OUT_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [1:0] O;
	assign O = I[25:24];
endmodule
module SB_T1_NORTH_SB_OUT_B1_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [2:0] O;
	assign O = I[29:27];
endmodule
module SB_T1_NORTH_SB_OUT_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [1:0] O;
	assign O = I[23:22];
endmodule
module SB_T1_NORTH_SB_OUT_B16_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [2:0] O;
	assign O = I[29:27];
endmodule
module SB_T1_NORTH_SB_OUT_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [1:0] O;
	assign O = I[23:22];
endmodule
module SB_T1_EAST_SB_OUT_B1_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [2:0] O;
	assign O = I[26:24];
endmodule
module SB_T1_EAST_SB_OUT_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [1:0] O;
	assign O = I[21:20];
endmodule
module SB_T1_EAST_SB_OUT_B16_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [2:0] O;
	assign O = I[26:24];
endmodule
module SB_T1_EAST_SB_OUT_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [1:0] O;
	assign O = I[21:20];
endmodule
module SB_T0_WEST_SB_OUT_B1_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [2:0] O;
	assign O = I[23:21];
endmodule
module SB_T0_WEST_SB_OUT_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [1:0] O;
	assign O = I[19:18];
endmodule
module SB_T0_WEST_SB_OUT_B16_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [2:0] O;
	assign O = I[23:21];
endmodule
module SB_T0_WEST_SB_OUT_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [1:0] O;
	assign O = I[19:18];
endmodule
module SB_T0_SOUTH_SB_OUT_B1_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [2:0] O;
	assign O = I[20:18];
endmodule
module SB_T0_SOUTH_SB_OUT_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [1:0] O;
	assign O = I[17:16];
endmodule
module SB_T0_SOUTH_SB_OUT_B16_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [2:0] O;
	assign O = I[20:18];
endmodule
module SB_T0_SOUTH_SB_OUT_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [1:0] O;
	assign O = I[17:16];
endmodule
module SB_T0_NORTH_SB_OUT_B1_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [2:0] O;
	assign O = I[17:15];
endmodule
module SB_T0_NORTH_SB_OUT_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [1:0] O;
	assign O = I[15:14];
endmodule
module SB_T0_NORTH_SB_OUT_B16_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [2:0] O;
	assign O = I[17:15];
endmodule
module SB_T0_NORTH_SB_OUT_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [1:0] O;
	assign O = I[15:14];
endmodule
module SB_T0_EAST_SB_OUT_B1_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [2:0] O;
	assign O = I[14:12];
endmodule
module SB_T0_EAST_SB_OUT_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [1:0] O;
	assign O = I[13:12];
endmodule
module SB_T0_EAST_SB_OUT_B16_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [2:0] O;
	assign O = I[14:12];
endmodule
module SB_T0_EAST_SB_OUT_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [1:0] O;
	assign O = I[13:12];
endmodule
module Register_unq9 (
	I,
	O,
	CE,
	CLK,
	ASYNCRESET
);
	input [10:0] I;
	output [10:0] O;
	input CE;
	input CLK;
	input ASYNCRESET;
	wire [10:0] reg_PR11_inst0__CE_out;
	regCE_arst #(
		.init(11'h000),
		.width(11)
	) reg_PR11_inst0__CE(
		.in(I),
		.ce(CE),
		.out(reg_PR11_inst0__CE_out),
		.clk(CLK),
		.arst(ASYNCRESET)
	);
	assign O = reg_PR11_inst0__CE_out;
endmodule
module Register_unq8 (
	I,
	O,
	CE,
	CLK,
	ASYNCRESET
);
	input [27:0] I;
	output [27:0] O;
	input CE;
	input CLK;
	input ASYNCRESET;
	wire [27:0] reg_PR28_inst0__CE_out;
	regCE_arst #(
		.init(28'h0000000),
		.width(28)
	) reg_PR28_inst0__CE(
		.in(I),
		.ce(CE),
		.out(reg_PR28_inst0__CE_out),
		.clk(CLK),
		.arst(ASYNCRESET)
	);
	assign O = reg_PR28_inst0__CE_out;
endmodule
module Register_unq7 (
	I,
	O,
	CE,
	CLK,
	ASYNCRESET
);
	input [24:0] I;
	output [24:0] O;
	input CE;
	input CLK;
	input ASYNCRESET;
	wire [24:0] reg_PR25_inst0__CE_out;
	regCE_arst #(
		.init(25'h0000000),
		.width(25)
	) reg_PR25_inst0__CE(
		.in(I),
		.ce(CE),
		.out(reg_PR25_inst0__CE_out),
		.clk(CLK),
		.arst(ASYNCRESET)
	);
	assign O = reg_PR25_inst0__CE_out;
endmodule
module Register_unq6 (
	I,
	O,
	CE,
	CLK,
	ASYNCRESET
);
	input [19:0] I;
	output [19:0] O;
	input CE;
	input CLK;
	input ASYNCRESET;
	wire [19:0] reg_PR20_inst0__CE_out;
	regCE_arst #(
		.init(20'h00000),
		.width(20)
	) reg_PR20_inst0__CE(
		.in(I),
		.ce(CE),
		.out(reg_PR20_inst0__CE_out),
		.clk(CLK),
		.arst(ASYNCRESET)
	);
	assign O = reg_PR20_inst0__CE_out;
endmodule
module Register_unq5 (
	I,
	O,
	CE,
	CLK,
	ASYNCRESET
);
	input [16:0] I;
	output [16:0] O;
	input CE;
	input CLK;
	input ASYNCRESET;
	wire [16:0] reg_PR17_inst0__CE_out;
	regCE_arst #(
		.init(17'h00000),
		.width(17)
	) reg_PR17_inst0__CE(
		.in(I),
		.ce(CE),
		.out(reg_PR17_inst0__CE_out),
		.clk(CLK),
		.arst(ASYNCRESET)
	);
	assign O = reg_PR17_inst0__CE_out;
endmodule
module Register_unq4 (
	I,
	O,
	CE,
	CLK,
	ASYNCRESET
);
	input [25:0] I;
	output [25:0] O;
	input CE;
	input CLK;
	input ASYNCRESET;
	wire [25:0] reg_PR26_inst0__CE_out;
	regCE_arst #(
		.init(26'h0000000),
		.width(26)
	) reg_PR26_inst0__CE(
		.in(I),
		.ce(CE),
		.out(reg_PR26_inst0__CE_out),
		.clk(CLK),
		.arst(ASYNCRESET)
	);
	assign O = reg_PR26_inst0__CE_out;
endmodule
module Register_unq3 (
	I,
	O,
	CE,
	CLK,
	ASYNCRESET
);
	input [31:0] I;
	output [31:0] O;
	input CE;
	input CLK;
	input ASYNCRESET;
	wire [31:0] reg_PR32_inst0__CE_out;
	regCE_arst #(
		.init(32'h00000000),
		.width(32)
	) reg_PR32_inst0__CE(
		.in(I),
		.ce(CE),
		.out(reg_PR32_inst0__CE_out),
		.clk(CLK),
		.arst(ASYNCRESET)
	);
	assign O = reg_PR32_inst0__CE_out;
endmodule
module Register_unq2 (
	value,
	O,
	en,
	CLK,
	ASYNCRESET
);
	input value;
	output O;
	input en;
	input CLK;
	input ASYNCRESET;
	wire [0:0] enable_mux$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] reg_PR1_inst0_out;
	coreir_mux #(.width(1)) enable_mux$coreir_commonlib_mux2x1_inst0$_join(
		.in0(reg_PR1_inst0_out[0]),
		.in1(value),
		.sel(en),
		.out(enable_mux$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_reg_arst #(
		.arst_posedge(1'b1),
		.clk_posedge(1'b1),
		.init(1'h0),
		.width(1)
	) reg_PR1_inst0(
		.clk(CLK),
		.arst(ASYNCRESET),
		.in(enable_mux$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.out(reg_PR1_inst0_out)
	);
	assign O = reg_PR1_inst0_out[0];
endmodule
module Register_unq11 (
	I,
	O,
	CE,
	CLK,
	ASYNCRESET
);
	input [17:0] I;
	output [17:0] O;
	input CE;
	input CLK;
	input ASYNCRESET;
	wire [17:0] reg_PR18_inst0__CE_out;
	regCE_arst #(
		.init(18'h00000),
		.width(18)
	) reg_PR18_inst0__CE(
		.in(I),
		.ce(CE),
		.out(reg_PR18_inst0__CE_out),
		.clk(CLK),
		.arst(ASYNCRESET)
	);
	assign O = reg_PR18_inst0__CE_out;
endmodule
module Register_unq10 (
	I,
	O,
	CE,
	CLK,
	ASYNCRESET
);
	input [29:0] I;
	output [29:0] O;
	input CE;
	input CLK;
	input ASYNCRESET;
	wire [29:0] reg_PR30_inst0__CE_out;
	regCE_arst #(
		.init(30'h00000000),
		.width(30)
	) reg_PR30_inst0__CE(
		.in(I),
		.ce(CE),
		.out(reg_PR30_inst0__CE_out),
		.clk(CLK),
		.arst(ASYNCRESET)
	);
	assign O = reg_PR30_inst0__CE_out;
endmodule
module Register_unq1 (
	value,
	O,
	en,
	CLK,
	ASYNCRESET
);
	input [15:0] value;
	output [15:0] O;
	input en;
	input CLK;
	input ASYNCRESET;
	wire [15:0] reg_PR16_inst0__CE_out;
	regCE_arst #(
		.init(16'h0000),
		.width(16)
	) reg_PR16_inst0__CE(
		.in(value),
		.ce(en),
		.out(reg_PR16_inst0__CE_out),
		.clk(CLK),
		.arst(ASYNCRESET)
	);
	assign O = reg_PR16_inst0__CE_out;
endmodule
module Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 (
	I,
	O,
	CLK,
	CE
);
	input [15:0] I;
	output [15:0] O;
	input CLK;
	input CE;
	wire [15:0] value__CE_out;
	regCE #(.width(16)) value__CE(
		.in(I),
		.ce(CE),
		.out(value__CE_out),
		.clk(CLK)
	);
	assign O = value__CE_out;
endmodule
module Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 (
	I,
	O,
	CLK,
	CE
);
	input [0:0] I;
	output [0:0] O;
	input CLK;
	input CE;
	wire [0:0] value__CE_out;
	regCE #(.width(1)) value__CE(
		.in(I),
		.ce(CE),
		.out(value__CE_out),
		.clk(CLK)
	);
	assign O = value__CE_out;
endmodule
module RegisterMode_unq1 (
	mode,
	const_,
	value,
	clk_en,
	config_we,
	config_data,
	O0,
	O1,
	CLK,
	ASYNCRESET
);
	input [1:0] mode;
	input const_;
	input value;
	input clk_en;
	input config_we;
	input config_data;
	output O0;
	output O1;
	input CLK;
	input ASYNCRESET;
	wire [0:0] Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out;
	wire Register_inst0_O;
	wire bit_const_0_None_out;
	wire bit_const_1_None_out;
	wire [1:0] const_0_2_out;
	wire [1:0] const_2_2_out;
	wire [1:0] const_3_2_out;
	wire magma_Bits_2_eq_inst0_out;
	wire magma_Bits_2_eq_inst1_out;
	wire magma_Bits_2_eq_inst2_out;
	coreir_mux #(.width(1)) Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(value),
		.in1(value),
		.sel(magma_Bits_2_eq_inst0_out),
		.out(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join(
		.in0(bit_const_0_None_out),
		.in1(clk_en),
		.sel(magma_Bits_2_eq_inst0_out),
		.out(Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(config_data),
		.sel(config_we),
		.out(Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_1_None_out),
		.sel(config_we),
		.out(Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Register_inst0_O),
		.in1(value),
		.sel(magma_Bits_2_eq_inst2_out),
		.out(Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst5$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Register_inst0_O),
		.in1(Register_inst0_O),
		.sel(magma_Bits_2_eq_inst2_out),
		.out(Mux2xBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst6$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(const_),
		.sel(magma_Bits_2_eq_inst1_out),
		.out(Mux2xBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst7$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(Register_inst0_O),
		.sel(magma_Bits_2_eq_inst1_out),
		.out(Mux2xBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	Register_unq2 Register_inst0(
		.value(Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.O(Register_inst0_O),
		.en(Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	corebit_const #(.value(1'b0)) bit_const_0_None(.out(bit_const_0_None_out));
	corebit_const #(.value(1'b1)) bit_const_1_None(.out(bit_const_1_None_out));
	coreir_const #(
		.value(2'h0),
		.width(2)
	) const_0_2(.out(const_0_2_out));
	coreir_const #(
		.value(2'h2),
		.width(2)
	) const_2_2(.out(const_2_2_out));
	coreir_const #(
		.value(2'h3),
		.width(2)
	) const_3_2(.out(const_3_2_out));
	coreir_eq #(.width(2)) magma_Bits_2_eq_inst0(
		.in0(mode),
		.in1(const_3_2_out),
		.out(magma_Bits_2_eq_inst0_out)
	);
	coreir_eq #(.width(2)) magma_Bits_2_eq_inst1(
		.in0(mode),
		.in1(const_0_2_out),
		.out(magma_Bits_2_eq_inst1_out)
	);
	coreir_eq #(.width(2)) magma_Bits_2_eq_inst2(
		.in0(mode),
		.in1(const_2_2_out),
		.out(magma_Bits_2_eq_inst2_out)
	);
	assign O0 = Mux2xBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out[0];
	assign O1 = Mux2xBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out[0];
endmodule
module RegisterMode (
	mode,
	const_,
	value,
	clk_en,
	config_we,
	config_data,
	O0,
	O1,
	CLK,
	ASYNCRESET
);
	input [1:0] mode;
	input [15:0] const_;
	input [15:0] value;
	input clk_en;
	input config_we;
	input [15:0] config_data;
	output [15:0] O0;
	output [15:0] O1;
	input CLK;
	input ASYNCRESET;
	wire [0:0] Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst5$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Register_inst0_O;
	wire bit_const_0_None_out;
	wire bit_const_1_None_out;
	wire [1:0] const_0_2_out;
	wire [1:0] const_2_2_out;
	wire [1:0] const_3_2_out;
	wire magma_Bits_2_eq_inst0_out;
	wire magma_Bits_2_eq_inst1_out;
	wire magma_Bits_2_eq_inst2_out;
	coreir_mux #(.width(1)) Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(bit_const_0_None_out),
		.in1(clk_en),
		.sel(magma_Bits_2_eq_inst0_out),
		.out(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_1_None_out),
		.sel(config_we),
		.out(Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(value),
		.in1(value),
		.sel(magma_Bits_2_eq_inst0_out),
		.out(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(config_data),
		.sel(config_we),
		.out(Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Register_inst0_O),
		.in1(value),
		.sel(magma_Bits_2_eq_inst2_out),
		.out(Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Register_inst0_O),
		.in1(Register_inst0_O),
		.sel(magma_Bits_2_eq_inst2_out),
		.out(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_),
		.sel(magma_Bits_2_eq_inst1_out),
		.out(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst5$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Register_inst0_O),
		.sel(magma_Bits_2_eq_inst1_out),
		.out(Mux2xBits16_inst5$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	Register_unq1 Register_inst0(
		.value(Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out),
		.O(Register_inst0_O),
		.en(Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	corebit_const #(.value(1'b0)) bit_const_0_None(.out(bit_const_0_None_out));
	corebit_const #(.value(1'b1)) bit_const_1_None(.out(bit_const_1_None_out));
	coreir_const #(
		.value(2'h0),
		.width(2)
	) const_0_2(.out(const_0_2_out));
	coreir_const #(
		.value(2'h2),
		.width(2)
	) const_2_2(.out(const_2_2_out));
	coreir_const #(
		.value(2'h3),
		.width(2)
	) const_3_2(.out(const_3_2_out));
	coreir_eq #(.width(2)) magma_Bits_2_eq_inst0(
		.in0(mode),
		.in1(const_3_2_out),
		.out(magma_Bits_2_eq_inst0_out)
	);
	coreir_eq #(.width(2)) magma_Bits_2_eq_inst1(
		.in0(mode),
		.in1(const_0_2_out),
		.out(magma_Bits_2_eq_inst1_out)
	);
	coreir_eq #(.width(2)) magma_Bits_2_eq_inst2(
		.in0(mode),
		.in1(const_2_2_out),
		.out(magma_Bits_2_eq_inst2_out)
	);
	assign O0 = Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out;
	assign O1 = Mux2xBits16_inst5$coreir_commonlib_mux2x16_inst0$_join_out;
endmodule
module Register (
	I,
	O,
	CE,
	CLK,
	ASYNCRESET
);
	input [3:0] I;
	output [3:0] O;
	input CE;
	input CLK;
	input ASYNCRESET;
	wire [3:0] reg_PR4_inst0__CE_out;
	regCE_arst #(
		.init(4'h0),
		.width(4)
	) reg_PR4_inst0__CE(
		.in(I),
		.ce(CE),
		.out(reg_PR4_inst0__CE_out),
		.clk(CLK),
		.arst(ASYNCRESET)
	);
	assign O = reg_PR4_inst0__CE_out;
endmodule
module RMUX_T2_WEST_B1_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[11];
endmodule
module RMUX_T2_WEST_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[11];
endmodule
module RMUX_T2_WEST_B16_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[11];
endmodule
module RMUX_T2_WEST_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[11];
endmodule
module RMUX_T2_SOUTH_B1_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[10];
endmodule
module RMUX_T2_SOUTH_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[10];
endmodule
module RMUX_T2_SOUTH_B16_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[10];
endmodule
module RMUX_T2_SOUTH_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[10];
endmodule
module RMUX_T2_NORTH_B1_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[9];
endmodule
module RMUX_T2_NORTH_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[9];
endmodule
module RMUX_T2_NORTH_B16_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[9];
endmodule
module RMUX_T2_NORTH_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[9];
endmodule
module RMUX_T2_EAST_B1_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[8];
endmodule
module RMUX_T2_EAST_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[8];
endmodule
module RMUX_T2_EAST_B16_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[8];
endmodule
module RMUX_T2_EAST_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[8];
endmodule
module RMUX_T1_WEST_B1_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[7];
endmodule
module RMUX_T1_WEST_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[7];
endmodule
module RMUX_T1_WEST_B16_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[7];
endmodule
module RMUX_T1_WEST_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[7];
endmodule
module RMUX_T1_SOUTH_B1_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[6];
endmodule
module RMUX_T1_SOUTH_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[6];
endmodule
module RMUX_T1_SOUTH_B16_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[6];
endmodule
module RMUX_T1_SOUTH_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[6];
endmodule
module RMUX_T1_NORTH_B1_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[5];
endmodule
module RMUX_T1_NORTH_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[5];
endmodule
module RMUX_T1_NORTH_B16_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[5];
endmodule
module RMUX_T1_NORTH_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[5];
endmodule
module RMUX_T1_EAST_B1_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[4];
endmodule
module RMUX_T1_EAST_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[4];
endmodule
module RMUX_T1_EAST_B16_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[4];
endmodule
module RMUX_T1_EAST_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[4];
endmodule
module RMUX_T0_WEST_B1_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[3];
endmodule
module RMUX_T0_WEST_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[3];
endmodule
module RMUX_T0_WEST_B16_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[3];
endmodule
module RMUX_T0_WEST_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[3];
endmodule
module RMUX_T0_SOUTH_B1_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[2];
endmodule
module RMUX_T0_SOUTH_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[2];
endmodule
module RMUX_T0_SOUTH_B16_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[2];
endmodule
module RMUX_T0_SOUTH_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[2];
endmodule
module RMUX_T0_NORTH_B1_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[1];
endmodule
module RMUX_T0_NORTH_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[1];
endmodule
module RMUX_T0_NORTH_B16_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[1];
endmodule
module RMUX_T0_NORTH_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[1];
endmodule
module RMUX_T0_EAST_B1_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[0];
endmodule
module RMUX_T0_EAST_B1_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[0];
endmodule
module RMUX_T0_EAST_B16_sel_unq1 (
	I,
	O
);
	input [29:0] I;
	output [0:0] O;
	assign O = I[0];
endmodule
module RMUX_T0_EAST_B16_sel (
	I,
	O
);
	input [31:0] I;
	output [0:0] O;
	assign O = I[0];
endmodule
module Or4x32 (
	I0,
	I1,
	I2,
	I3,
	O
);
	input [31:0] I0;
	input [31:0] I1;
	input [31:0] I2;
	input [31:0] I3;
	output [31:0] O;
	wire orr_inst0_out;
	wire orr_inst1_out;
	wire orr_inst10_out;
	wire orr_inst11_out;
	wire orr_inst12_out;
	wire orr_inst13_out;
	wire orr_inst14_out;
	wire orr_inst15_out;
	wire orr_inst16_out;
	wire orr_inst17_out;
	wire orr_inst18_out;
	wire orr_inst19_out;
	wire orr_inst2_out;
	wire orr_inst20_out;
	wire orr_inst21_out;
	wire orr_inst22_out;
	wire orr_inst23_out;
	wire orr_inst24_out;
	wire orr_inst25_out;
	wire orr_inst26_out;
	wire orr_inst27_out;
	wire orr_inst28_out;
	wire orr_inst29_out;
	wire orr_inst3_out;
	wire orr_inst30_out;
	wire orr_inst31_out;
	wire orr_inst4_out;
	wire orr_inst5_out;
	wire orr_inst6_out;
	wire orr_inst7_out;
	wire orr_inst8_out;
	wire orr_inst9_out;
	wire [3:0] orr_inst0_in;
	assign orr_inst0_in = {I3[0], I2[0], I1[0], I0[0]};
	coreir_orr #(.width(4)) orr_inst0(
		.in(orr_inst0_in),
		.out(orr_inst0_out)
	);
	wire [3:0] orr_inst1_in;
	assign orr_inst1_in = {I3[1], I2[1], I1[1], I0[1]};
	coreir_orr #(.width(4)) orr_inst1(
		.in(orr_inst1_in),
		.out(orr_inst1_out)
	);
	wire [3:0] orr_inst10_in;
	assign orr_inst10_in = {I3[10], I2[10], I1[10], I0[10]};
	coreir_orr #(.width(4)) orr_inst10(
		.in(orr_inst10_in),
		.out(orr_inst10_out)
	);
	wire [3:0] orr_inst11_in;
	assign orr_inst11_in = {I3[11], I2[11], I1[11], I0[11]};
	coreir_orr #(.width(4)) orr_inst11(
		.in(orr_inst11_in),
		.out(orr_inst11_out)
	);
	wire [3:0] orr_inst12_in;
	assign orr_inst12_in = {I3[12], I2[12], I1[12], I0[12]};
	coreir_orr #(.width(4)) orr_inst12(
		.in(orr_inst12_in),
		.out(orr_inst12_out)
	);
	wire [3:0] orr_inst13_in;
	assign orr_inst13_in = {I3[13], I2[13], I1[13], I0[13]};
	coreir_orr #(.width(4)) orr_inst13(
		.in(orr_inst13_in),
		.out(orr_inst13_out)
	);
	wire [3:0] orr_inst14_in;
	assign orr_inst14_in = {I3[14], I2[14], I1[14], I0[14]};
	coreir_orr #(.width(4)) orr_inst14(
		.in(orr_inst14_in),
		.out(orr_inst14_out)
	);
	wire [3:0] orr_inst15_in;
	assign orr_inst15_in = {I3[15], I2[15], I1[15], I0[15]};
	coreir_orr #(.width(4)) orr_inst15(
		.in(orr_inst15_in),
		.out(orr_inst15_out)
	);
	wire [3:0] orr_inst16_in;
	assign orr_inst16_in = {I3[16], I2[16], I1[16], I0[16]};
	coreir_orr #(.width(4)) orr_inst16(
		.in(orr_inst16_in),
		.out(orr_inst16_out)
	);
	wire [3:0] orr_inst17_in;
	assign orr_inst17_in = {I3[17], I2[17], I1[17], I0[17]};
	coreir_orr #(.width(4)) orr_inst17(
		.in(orr_inst17_in),
		.out(orr_inst17_out)
	);
	wire [3:0] orr_inst18_in;
	assign orr_inst18_in = {I3[18], I2[18], I1[18], I0[18]};
	coreir_orr #(.width(4)) orr_inst18(
		.in(orr_inst18_in),
		.out(orr_inst18_out)
	);
	wire [3:0] orr_inst19_in;
	assign orr_inst19_in = {I3[19], I2[19], I1[19], I0[19]};
	coreir_orr #(.width(4)) orr_inst19(
		.in(orr_inst19_in),
		.out(orr_inst19_out)
	);
	wire [3:0] orr_inst2_in;
	assign orr_inst2_in = {I3[2], I2[2], I1[2], I0[2]};
	coreir_orr #(.width(4)) orr_inst2(
		.in(orr_inst2_in),
		.out(orr_inst2_out)
	);
	wire [3:0] orr_inst20_in;
	assign orr_inst20_in = {I3[20], I2[20], I1[20], I0[20]};
	coreir_orr #(.width(4)) orr_inst20(
		.in(orr_inst20_in),
		.out(orr_inst20_out)
	);
	wire [3:0] orr_inst21_in;
	assign orr_inst21_in = {I3[21], I2[21], I1[21], I0[21]};
	coreir_orr #(.width(4)) orr_inst21(
		.in(orr_inst21_in),
		.out(orr_inst21_out)
	);
	wire [3:0] orr_inst22_in;
	assign orr_inst22_in = {I3[22], I2[22], I1[22], I0[22]};
	coreir_orr #(.width(4)) orr_inst22(
		.in(orr_inst22_in),
		.out(orr_inst22_out)
	);
	wire [3:0] orr_inst23_in;
	assign orr_inst23_in = {I3[23], I2[23], I1[23], I0[23]};
	coreir_orr #(.width(4)) orr_inst23(
		.in(orr_inst23_in),
		.out(orr_inst23_out)
	);
	wire [3:0] orr_inst24_in;
	assign orr_inst24_in = {I3[24], I2[24], I1[24], I0[24]};
	coreir_orr #(.width(4)) orr_inst24(
		.in(orr_inst24_in),
		.out(orr_inst24_out)
	);
	wire [3:0] orr_inst25_in;
	assign orr_inst25_in = {I3[25], I2[25], I1[25], I0[25]};
	coreir_orr #(.width(4)) orr_inst25(
		.in(orr_inst25_in),
		.out(orr_inst25_out)
	);
	wire [3:0] orr_inst26_in;
	assign orr_inst26_in = {I3[26], I2[26], I1[26], I0[26]};
	coreir_orr #(.width(4)) orr_inst26(
		.in(orr_inst26_in),
		.out(orr_inst26_out)
	);
	wire [3:0] orr_inst27_in;
	assign orr_inst27_in = {I3[27], I2[27], I1[27], I0[27]};
	coreir_orr #(.width(4)) orr_inst27(
		.in(orr_inst27_in),
		.out(orr_inst27_out)
	);
	wire [3:0] orr_inst28_in;
	assign orr_inst28_in = {I3[28], I2[28], I1[28], I0[28]};
	coreir_orr #(.width(4)) orr_inst28(
		.in(orr_inst28_in),
		.out(orr_inst28_out)
	);
	wire [3:0] orr_inst29_in;
	assign orr_inst29_in = {I3[29], I2[29], I1[29], I0[29]};
	coreir_orr #(.width(4)) orr_inst29(
		.in(orr_inst29_in),
		.out(orr_inst29_out)
	);
	wire [3:0] orr_inst3_in;
	assign orr_inst3_in = {I3[3], I2[3], I1[3], I0[3]};
	coreir_orr #(.width(4)) orr_inst3(
		.in(orr_inst3_in),
		.out(orr_inst3_out)
	);
	wire [3:0] orr_inst30_in;
	assign orr_inst30_in = {I3[30], I2[30], I1[30], I0[30]};
	coreir_orr #(.width(4)) orr_inst30(
		.in(orr_inst30_in),
		.out(orr_inst30_out)
	);
	wire [3:0] orr_inst31_in;
	assign orr_inst31_in = {I3[31], I2[31], I1[31], I0[31]};
	coreir_orr #(.width(4)) orr_inst31(
		.in(orr_inst31_in),
		.out(orr_inst31_out)
	);
	wire [3:0] orr_inst4_in;
	assign orr_inst4_in = {I3[4], I2[4], I1[4], I0[4]};
	coreir_orr #(.width(4)) orr_inst4(
		.in(orr_inst4_in),
		.out(orr_inst4_out)
	);
	wire [3:0] orr_inst5_in;
	assign orr_inst5_in = {I3[5], I2[5], I1[5], I0[5]};
	coreir_orr #(.width(4)) orr_inst5(
		.in(orr_inst5_in),
		.out(orr_inst5_out)
	);
	wire [3:0] orr_inst6_in;
	assign orr_inst6_in = {I3[6], I2[6], I1[6], I0[6]};
	coreir_orr #(.width(4)) orr_inst6(
		.in(orr_inst6_in),
		.out(orr_inst6_out)
	);
	wire [3:0] orr_inst7_in;
	assign orr_inst7_in = {I3[7], I2[7], I1[7], I0[7]};
	coreir_orr #(.width(4)) orr_inst7(
		.in(orr_inst7_in),
		.out(orr_inst7_out)
	);
	wire [3:0] orr_inst8_in;
	assign orr_inst8_in = {I3[8], I2[8], I1[8], I0[8]};
	coreir_orr #(.width(4)) orr_inst8(
		.in(orr_inst8_in),
		.out(orr_inst8_out)
	);
	wire [3:0] orr_inst9_in;
	assign orr_inst9_in = {I3[9], I2[9], I1[9], I0[9]};
	coreir_orr #(.width(4)) orr_inst9(
		.in(orr_inst9_in),
		.out(orr_inst9_out)
	);
	assign O = {orr_inst31_out, orr_inst30_out, orr_inst29_out, orr_inst28_out, orr_inst27_out, orr_inst26_out, orr_inst25_out, orr_inst24_out, orr_inst23_out, orr_inst22_out, orr_inst21_out, orr_inst20_out, orr_inst19_out, orr_inst18_out, orr_inst17_out, orr_inst16_out, orr_inst15_out, orr_inst14_out, orr_inst13_out, orr_inst12_out, orr_inst11_out, orr_inst10_out, orr_inst9_out, orr_inst8_out, orr_inst7_out, orr_inst6_out, orr_inst5_out, orr_inst4_out, orr_inst3_out, orr_inst2_out, orr_inst1_out, orr_inst0_out};
endmodule
module MuxWrapper_1_16 (
	I,
	O
);
	input [15:0] I;
	output [15:0] O;
	assign O = I;
endmodule
module MuxWrapper_1_1 (
	I,
	O
);
	input [0:0] I;
	output [0:0] O;
	assign O = I;
endmodule
module Tile_io_core (
	tile_id,
	glb2io_1,
	f2io_1,
	io2glb_1,
	io2f_1,
	glb2io_16,
	f2io_16,
	io2glb_16,
	io2f_16,
	hi,
	lo
);
	input [15:0] tile_id;
	input [0:0] glb2io_1;
	input [0:0] f2io_1;
	output [0:0] io2glb_1;
	output [0:0] io2f_1;
	input [15:0] glb2io_16;
	input [15:0] f2io_16;
	output [15:0] io2glb_16;
	output [15:0] io2f_16;
	output [8:0] hi;
	output [7:0] lo;
	wire [0:0] CB_f2io_1$WIRE_CB_f2io_1_O;
	wire [15:0] CB_f2io_16$WIRE_CB_f2io_16_O;
	wire [7:0] const_0_8_out;
	wire [8:0] const_511_9_out;
	wire [15:0] io_core_inst0_io2glb_16;
	wire [0:0] io_core_inst0_io2glb_1;
	wire [15:0] io_core_inst0_io2f_16;
	wire [0:0] io_core_inst0_io2f_1;
	MuxWrapper_1_1 CB_f2io_1$WIRE_CB_f2io_1(
		.I(f2io_1),
		.O(CB_f2io_1$WIRE_CB_f2io_1_O)
	);
	MuxWrapper_1_16 CB_f2io_16$WIRE_CB_f2io_16(
		.I(f2io_16),
		.O(CB_f2io_16$WIRE_CB_f2io_16_O)
	);
	coreir_const #(
		.value(8'h00),
		.width(8)
	) const_0_8(.out(const_0_8_out));
	coreir_const #(
		.value(9'h1ff),
		.width(9)
	) const_511_9(.out(const_511_9_out));
	io_core io_core_inst0(
		.glb2io_16(glb2io_16),
		.glb2io_1(glb2io_1),
		.io2glb_16(io_core_inst0_io2glb_16),
		.io2glb_1(io_core_inst0_io2glb_1),
		.f2io_16(CB_f2io_16$WIRE_CB_f2io_16_O),
		.f2io_1(CB_f2io_1$WIRE_CB_f2io_1_O),
		.io2f_16(io_core_inst0_io2f_16),
		.io2f_1(io_core_inst0_io2f_1)
	);
	assign io2glb_1 = io_core_inst0_io2glb_1;
	assign io2f_1 = io_core_inst0_io2f_1;
	assign io2glb_16 = io_core_inst0_io2glb_16;
	assign io2f_16 = io_core_inst0_io2f_16;
	assign hi = const_511_9_out;
	assign lo = const_0_8_out;
endmodule
module MuxWithDefaultWrapper_8_32_8_0 (
	EN,
	I_0,
	I_1,
	I_2,
	I_3,
	I_4,
	I_5,
	I_6,
	I_7,
	O,
	S
);
	input [0:0] EN;
	input [31:0] I_0;
	input [31:0] I_1;
	input [31:0] I_2;
	input [31:0] I_3;
	input [31:0] I_4;
	input [31:0] I_5;
	input [31:0] I_6;
	input [31:0] I_7;
	output [31:0] O;
	input [7:0] S;
	wire [31:0] MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
	wire [31:0] MuxWrapper_8_32_inst0$Mux8xBits32_inst0$coreir_commonlib_mux8x32_inst0_out;
	wire [2:0] MuxWrapper_8_32_inst0_S_in;
	wire [31:0] const_0_32_out;
	wire [7:0] const_8_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_ult_inst0_out;
	wire [7:0] self_S_out;
	coreir_mux #(.width(32)) MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join(
		.in0(const_0_32_out),
		.in1(MuxWrapper_8_32_inst0$Mux8xBits32_inst0$coreir_commonlib_mux8x32_inst0_out),
		.sel(magma_Bit_and_inst0_out),
		.out(MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out)
	);
	commonlib_muxn__N8__width32 MuxWrapper_8_32_inst0$Mux8xBits32_inst0$coreir_commonlib_mux8x32_inst0(
		.in_data_0(I_0),
		.in_data_1(I_1),
		.in_data_2(I_2),
		.in_data_3(I_3),
		.in_data_4(I_4),
		.in_data_5(I_5),
		.in_data_6(I_6),
		.in_data_7(I_7),
		.in_sel(MuxWrapper_8_32_inst0_S_in),
		.out(MuxWrapper_8_32_inst0$Mux8xBits32_inst0$coreir_commonlib_mux8x32_inst0_out)
	);
	mantle_wire__typeBitIn3 MuxWrapper_8_32_inst0_S(
		.in(MuxWrapper_8_32_inst0_S_in),
		.out(self_S_out[2:0])
	);
	coreir_const #(
		.value(32'h00000000),
		.width(32)
	) const_0_32(.out(const_0_32_out));
	coreir_const #(
		.value(8'h08),
		.width(8)
	) const_8_8(.out(const_8_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_ult_inst0_out),
		.in1(EN[0]),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_ult #(.width(8)) magma_Bits_8_ult_inst0(
		.in0(S),
		.in1(const_8_8_out),
		.out(magma_Bits_8_ult_inst0_out)
	);
	mantle_wire__typeBit8 self_S(
		.in(S),
		.out(self_S_out)
	);
	assign O = MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
endmodule
module MuxWithDefaultWrapper_11_32_8_0 (
	EN,
	I_0,
	I_1,
	I_10,
	I_2,
	I_3,
	I_4,
	I_5,
	I_6,
	I_7,
	I_8,
	I_9,
	O,
	S
);
	input [0:0] EN;
	input [31:0] I_0;
	input [31:0] I_1;
	input [31:0] I_10;
	input [31:0] I_2;
	input [31:0] I_3;
	input [31:0] I_4;
	input [31:0] I_5;
	input [31:0] I_6;
	input [31:0] I_7;
	input [31:0] I_8;
	input [31:0] I_9;
	output [31:0] O;
	input [7:0] S;
	wire [31:0] MuxWrapper_11_32_inst0$Mux11xBits32_inst0$coreir_commonlib_mux11x32_inst0_out;
	wire [3:0] MuxWrapper_11_32_inst0_S_in;
	wire [31:0] MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
	wire [31:0] const_0_32_out;
	wire [7:0] const_11_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_ult_inst0_out;
	wire [7:0] self_S_out;
	commonlib_muxn__N11__width32 MuxWrapper_11_32_inst0$Mux11xBits32_inst0$coreir_commonlib_mux11x32_inst0(
		.in_data_0(I_0),
		.in_data_1(I_1),
		.in_data_10(I_10),
		.in_data_2(I_2),
		.in_data_3(I_3),
		.in_data_4(I_4),
		.in_data_5(I_5),
		.in_data_6(I_6),
		.in_data_7(I_7),
		.in_data_8(I_8),
		.in_data_9(I_9),
		.in_sel(MuxWrapper_11_32_inst0_S_in),
		.out(MuxWrapper_11_32_inst0$Mux11xBits32_inst0$coreir_commonlib_mux11x32_inst0_out)
	);
	mantle_wire__typeBitIn4 MuxWrapper_11_32_inst0_S(
		.in(MuxWrapper_11_32_inst0_S_in),
		.out(self_S_out[3:0])
	);
	coreir_mux #(.width(32)) MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join(
		.in0(const_0_32_out),
		.in1(MuxWrapper_11_32_inst0$Mux11xBits32_inst0$coreir_commonlib_mux11x32_inst0_out),
		.sel(magma_Bit_and_inst0_out),
		.out(MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out)
	);
	coreir_const #(
		.value(32'h00000000),
		.width(32)
	) const_0_32(.out(const_0_32_out));
	coreir_const #(
		.value(8'h0b),
		.width(8)
	) const_11_8(.out(const_11_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_ult_inst0_out),
		.in1(EN[0]),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_ult #(.width(8)) magma_Bits_8_ult_inst0(
		.in0(S),
		.in1(const_11_8_out),
		.out(magma_Bits_8_ult_inst0_out)
	);
	mantle_wire__typeBit8 self_S(
		.in(S),
		.out(self_S_out)
	);
	assign O = MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
endmodule
module Chain (
	accessor_output,
	chain_data_in,
	chain_en,
	clk_en,
	curr_tile_data_out,
	flush,
	data_out_tile
);
	input wire [1:0] accessor_output;
	input wire [31:0] chain_data_in;
	input wire chain_en;
	input wire clk_en;
	input wire [31:0] curr_tile_data_out;
	input wire flush;
	output reg [31:0] data_out_tile;
	always @(*) begin
		if (accessor_output[0])
			data_out_tile[0+:16] = curr_tile_data_out[0+:16];
		else if (chain_en)
			data_out_tile[0+:16] = chain_data_in[0+:16];
		else
			data_out_tile[0+:16] = 16'h0000;
		if (accessor_output[1])
			data_out_tile[16+:16] = curr_tile_data_out[16+:16];
		else if (chain_en)
			data_out_tile[16+:16] = chain_data_in[16+:16];
		else
			data_out_tile[16+:16] = 16'h0000;
	end
endmodule
module LakeTop (
	clk,
	clk_en,
	config_addr_in,
	config_data_in,
	config_en,
	config_read,
	config_write,
	flush,
	input_width_16_num_0,
	input_width_16_num_1,
	input_width_16_num_2,
	input_width_16_num_3,
	input_width_1_num_0,
	input_width_1_num_1,
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality,
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges,
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable,
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr,
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides,
	mode,
	rst_n,
	tile_en,
	config_data_out,
	output_width_16_num_0,
	output_width_16_num_1,
	output_width_1_num_0,
	output_width_1_num_1,
	output_width_1_num_2
);
	input wire clk;
	input wire clk_en;
	input wire [7:0] config_addr_in;
	input wire [31:0] config_data_in;
	input wire config_en;
	input wire config_read;
	input wire config_write;
	input wire flush;
	input wire [15:0] input_width_16_num_0;
	input wire [15:0] input_width_16_num_1;
	input wire [15:0] input_width_16_num_2;
	input wire [15:0] input_width_16_num_3;
	input wire input_width_1_num_0;
	input wire input_width_1_num_1;
	input wire [3:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality;
	input wire [95:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges;
	input wire mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable;
	input wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr;
	input wire [95:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr;
	input wire [23:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr;
	input wire [23:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr;
	input wire [23:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr;
	input wire [23:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides;
	input wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr;
	input wire [95:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides;
	input wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr;
	input wire [95:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality;
	input wire [95:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality;
	input wire [95:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges;
	input wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr;
	input wire [95:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides;
	input wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr;
	input wire [95:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality;
	input wire [95:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality;
	input wire [95:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges;
	input wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr;
	input wire [47:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr;
	input wire [47:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr;
	input wire [47:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr;
	input wire [47:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality;
	// input wire [95:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality;
	// input wire [95:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges;
	// input wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr;
	// input wire [95:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides;
	// input wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr;
	// input wire [95:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality;
	// input wire [95:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality;
	// input wire [95:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr;
	// input wire [23:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr;
	// input wire [23:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides;
	// input wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr;
	// input wire [95:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides;
	// input wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr;
	// input wire [95:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr;
	// input wire [23:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr;
	// input wire [23:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides;
	input wire [1:0] mode;
	input wire rst_n;
	input wire tile_en;
	output wire [31:0] config_data_out;
	output reg [15:0] output_width_16_num_0;
	output reg [15:0] output_width_16_num_1;
	output reg output_width_1_num_0;
	output reg output_width_1_num_1;
	output reg output_width_1_num_2;
	wire [15:0] config_data_in_shrt;
	wire [15:0] config_data_out_shrt;
	wire [7:0] config_seq_addr_out;
	wire config_seq_clk;
	wire config_seq_clk_en;
	reg [31:0] config_seq_rd_data_stg;
	wire config_seq_ren_out;
	wire config_seq_wen_out;
	wire [31:0] config_seq_wr_data;
	wire gclk;
	wire mem_ctrl_stencil_valid_flat_clk;
	wire mem_ctrl_stencil_valid_flat_stencil_valid_f_;
	wire [7:0] mem_ctrl_strg_ram_flat_addr_out_lifted;
	wire mem_ctrl_strg_ram_flat_clk;
	reg [31:0] mem_ctrl_strg_ram_flat_data_from_strg_lifted;
	wire [15:0] mem_ctrl_strg_ram_flat_data_out_f_;
	wire [31:0] mem_ctrl_strg_ram_flat_data_to_strg_lifted;
	wire mem_ctrl_strg_ram_flat_ready_f_;
	wire mem_ctrl_strg_ram_flat_ren_to_strg_lifted;
	wire mem_ctrl_strg_ram_flat_valid_out_f_;
	wire mem_ctrl_strg_ram_flat_wen_to_strg_lifted;
	wire mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_0;
	wire mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_1;
	wire mem_ctrl_strg_ub_vec_flat_clk;
	reg [31:0] mem_ctrl_strg_ub_vec_flat_data_from_strg_lifted;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_data_out_f_0;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_data_out_f_1;
	wire [31:0] mem_ctrl_strg_ub_vec_flat_data_to_strg_lifted;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_rd_addr_out_lifted;
	wire mem_ctrl_strg_ub_vec_flat_ren_to_strg_lifted;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_tmp0_rdaddr_lifted;
	wire mem_ctrl_strg_ub_vec_flat_tmp0_rden_lifted;
	wire mem_ctrl_strg_ub_vec_flat_wen_to_strg_lifted;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_wr_addr_out_lifted;
	wire memory_0_clk;
	wire memory_0_clk_en;
	reg [31:0] memory_0_data_in_p0;
	wire [31:0] memory_0_data_out_p0;
	wire [31:0] memory_0_data_out_p1;
	reg [7:0] memory_0_read_addr_p0;
	reg [7:0] memory_0_read_addr_p1;
	reg memory_0_read_enable_p0;
	reg memory_0_read_enable_p1;
	reg [7:0] memory_0_write_addr_p0;
	reg memory_0_write_enable_p0;
	assign gclk = clk & tile_en;
	assign mem_ctrl_strg_ub_vec_flat_clk = gclk & (mode == 2'h0);
	assign mem_ctrl_strg_ram_flat_clk = gclk & (mode == 2'h1);
	assign mem_ctrl_stencil_valid_flat_clk = gclk;
	always @(*) begin
		output_width_1_num_0 = 1'h0;
		if (mode == 2'h0)
			output_width_1_num_0 = mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_0;
		else if (mode == 2'h1)
			output_width_1_num_0 = mem_ctrl_strg_ram_flat_ready_f_;
	end
	always @(*) begin
		output_width_1_num_1 = 1'h0;
		if (mode == 2'h0)
			output_width_1_num_1 = mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_1;
		else if (mode == 2'h1)
			output_width_1_num_1 = mem_ctrl_strg_ram_flat_valid_out_f_;
	end
	always @(*) begin
		output_width_1_num_2 = 1'h0;
		output_width_1_num_2 = mem_ctrl_stencil_valid_flat_stencil_valid_f_;
	end
	always @(*) begin
		output_width_16_num_0 = 16'h0000;
		if (mode == 2'h0)
			output_width_16_num_0 = mem_ctrl_strg_ub_vec_flat_data_out_f_0;
		else if (mode == 2'h1)
			output_width_16_num_0 = mem_ctrl_strg_ram_flat_data_out_f_;
	end
	always @(*) begin
		output_width_16_num_1 = 16'h0000;
		output_width_16_num_1 = mem_ctrl_strg_ub_vec_flat_data_out_f_1;
	end
	assign memory_0_clk = gclk;
	always @(*) begin
		memory_0_data_in_p0 = 32'h00000000;
		memory_0_write_addr_p0 = 8'h00;
		memory_0_write_enable_p0 = 1'h0;
		memory_0_read_addr_p0 = 8'h00;
		memory_0_read_enable_p0 = 1'h0;
		if (|config_en) begin
			memory_0_data_in_p0 = config_seq_wr_data;
			memory_0_write_addr_p0 = config_seq_addr_out;
			memory_0_write_enable_p0 = config_seq_wen_out;
			memory_0_read_addr_p0 = config_seq_addr_out;
			memory_0_read_enable_p0 = config_seq_ren_out;
		end
		else if (mode == 2'h0) begin
			memory_0_data_in_p0 = mem_ctrl_strg_ub_vec_flat_data_to_strg_lifted;
			memory_0_write_addr_p0 = mem_ctrl_strg_ub_vec_flat_wr_addr_out_lifted;
			memory_0_write_enable_p0 = mem_ctrl_strg_ub_vec_flat_wen_to_strg_lifted;
			memory_0_read_addr_p0 = mem_ctrl_strg_ub_vec_flat_tmp0_rdaddr_lifted;
			memory_0_read_enable_p0 = mem_ctrl_strg_ub_vec_flat_tmp0_rden_lifted;
		end
		else if (mode == 2'h1) begin
			memory_0_data_in_p0 = mem_ctrl_strg_ram_flat_data_to_strg_lifted;
			memory_0_write_addr_p0 = mem_ctrl_strg_ram_flat_addr_out_lifted;
			memory_0_write_enable_p0 = mem_ctrl_strg_ram_flat_wen_to_strg_lifted;
			memory_0_read_addr_p0 = mem_ctrl_strg_ram_flat_addr_out_lifted;
			memory_0_read_enable_p0 = mem_ctrl_strg_ram_flat_ren_to_strg_lifted;
		end
	end
	always @(*) begin
		mem_ctrl_strg_ram_flat_data_from_strg_lifted = memory_0_data_out_p0;
		config_seq_rd_data_stg = memory_0_data_out_p0;
	end
	always @(*) begin
		memory_0_read_addr_p1 = 8'h00;
		memory_0_read_enable_p1 = 1'h0;
		if (mode == 2'h0) begin
			memory_0_read_addr_p1 = mem_ctrl_strg_ub_vec_flat_rd_addr_out_lifted;
			memory_0_read_enable_p1 = mem_ctrl_strg_ub_vec_flat_ren_to_strg_lifted;
		end
	end
	always @(*) mem_ctrl_strg_ub_vec_flat_data_from_strg_lifted = memory_0_data_out_p1;
	assign config_data_in_shrt = config_data_in[15:0];
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	assign config_data_out[0+:32] = sv2v_cast_32(config_data_out_shrt[0+:16]);
	assign config_seq_clk = gclk;
	assign config_seq_clk_en = clk_en | |config_en;
	assign memory_0_clk_en = clk_en | |config_en;
	strg_ub_vec_flat mem_ctrl_strg_ub_vec_flat(
		.chain_data_in_f_0(input_width_16_num_0),
		.chain_data_in_f_1(input_width_16_num_1),
		.clk(mem_ctrl_strg_ub_vec_flat_clk),
		.clk_en(clk_en),
		.data_from_strg_lifted(mem_ctrl_strg_ub_vec_flat_data_from_strg_lifted),
		.data_in_f_0(input_width_16_num_2),
		.data_in_f_1(input_width_16_num_3),
		.flush(flush),
		.rst_n(rst_n),
		.strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr),
		.strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides),
		.strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr),
		.strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides),
		.strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr),
		.strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides),
		.strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr),
		.strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides),
		.strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable),
		.strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr),
		.strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides),
		.strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable),
		.strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr),
		.strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides),
		.strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality),
		.strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges),
		.strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality),
		.strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges),
		.strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable),
		.strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr),
		.strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides),
		.strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable),
		.strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr),
		.strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides),
		.strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality),
		.strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges),
		.strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality),
		.strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges),
		.strg_ub_vec_inst_chain_chain_en(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en),
		.strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr),
		.strg_ub_vec_inst_sram_only_input_addr_gen_0_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides),
		.strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr),
		.strg_ub_vec_inst_sram_only_input_addr_gen_1_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides),
		.strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr),
		.strg_ub_vec_inst_sram_only_output_addr_gen_0_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides),
		.strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr),
		.strg_ub_vec_inst_sram_only_output_addr_gen_1_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides),
		// .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality),
		// .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges),
		// .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality),
		// .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges),
		// .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable),
		// .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr),
		// .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides),
		// .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable),
		// .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr),
		// .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides),
		// .strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality),
		// .strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges),
		// .strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality),
		// .strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges),
		// .strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr),
		// .strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides),
		// .strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr),
		// .strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides),
		// .strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable),
		// .strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr),
		// .strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides),
		// .strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable),
		// .strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr),
		// .strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides),
		// .strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr),
		// .strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides),
		// .strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr),
		// .strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides),
		.accessor_output_f_b_0(mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_0),
		.accessor_output_f_b_1(mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_1),
		.data_out_f_0(mem_ctrl_strg_ub_vec_flat_data_out_f_0),
		.data_out_f_1(mem_ctrl_strg_ub_vec_flat_data_out_f_1),
		.data_to_strg_lifted(mem_ctrl_strg_ub_vec_flat_data_to_strg_lifted),
		.rd_addr_out_lifted(mem_ctrl_strg_ub_vec_flat_rd_addr_out_lifted),
		.ren_to_strg_lifted(mem_ctrl_strg_ub_vec_flat_ren_to_strg_lifted),
		.tmp0_rdaddr_lifted(mem_ctrl_strg_ub_vec_flat_tmp0_rdaddr_lifted),
		.tmp0_rden_lifted(mem_ctrl_strg_ub_vec_flat_tmp0_rden_lifted),
		.wen_to_strg_lifted(mem_ctrl_strg_ub_vec_flat_wen_to_strg_lifted),
		.wr_addr_out_lifted(mem_ctrl_strg_ub_vec_flat_wr_addr_out_lifted)
	);
	strg_ram_flat mem_ctrl_strg_ram_flat(
		.clk(mem_ctrl_strg_ram_flat_clk),
		.clk_en(clk_en),
		.data_from_strg_lifted(mem_ctrl_strg_ram_flat_data_from_strg_lifted),
		.data_in_f_(input_width_16_num_0),
		.flush(flush),
		.rd_addr_in_f_(input_width_16_num_1),
		.ren_f_(input_width_1_num_0),
		.rst_n(rst_n),
		.wen_f_(input_width_1_num_1),
		.wr_addr_in_f_(input_width_16_num_2),
		.addr_out_lifted(mem_ctrl_strg_ram_flat_addr_out_lifted),
		.data_out_f_(mem_ctrl_strg_ram_flat_data_out_f_),
		.data_to_strg_lifted(mem_ctrl_strg_ram_flat_data_to_strg_lifted),
		.ready_f_(mem_ctrl_strg_ram_flat_ready_f_),
		.ren_to_strg_lifted(mem_ctrl_strg_ram_flat_ren_to_strg_lifted),
		.valid_out_f_(mem_ctrl_strg_ram_flat_valid_out_f_),
		.wen_to_strg_lifted(mem_ctrl_strg_ram_flat_wen_to_strg_lifted)
	);
	stencil_valid_flat mem_ctrl_stencil_valid_flat(
		.clk(mem_ctrl_stencil_valid_flat_clk),
		.clk_en(clk_en),
		.flush(flush),
		.rst_n(rst_n),
		.stencil_valid_inst_loops_stencil_valid_dimensionality(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality),
		.stencil_valid_inst_loops_stencil_valid_ranges(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges),
		.stencil_valid_inst_stencil_valid_sched_gen_enable(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable),
		.stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr),
		.stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides),
		.stencil_valid_f_(mem_ctrl_stencil_valid_flat_stencil_valid_f_)
	);
	sky130_sram_1kbyte_1rw1r_32x256_8 memory_0(
		.clk0(memory_0_clk),
		.csb0(~memory_0_clk_en),
		.web0(~memory_0_write_enable_p0),
		.wmask0(4'b1111),
		.addr0((memory_0_write_enable_p0 ? memory_0_write_addr_p0 : memory_0_read_addr_p0)),
		.din0(memory_0_data_in_p0),
		.dout0(memory_0_data_out_p0),
		.clk1(memory_0_clk),
		.csb1(~memory_0_clk_en),
		.addr1(memory_0_read_addr_p1),
		.dout1(memory_0_data_out_p1)
	);
	storage_config_seq config_seq(
		.clk(config_seq_clk),
		.clk_en(config_seq_clk_en),
		.config_addr_in(config_addr_in),
		.config_data_in(config_data_in_shrt),
		.config_en(config_en),
		.config_rd(config_read),
		.config_wr(config_write),
		.flush(flush),
		.rd_data_stg(config_seq_rd_data_stg),
		.rst_n(rst_n),
		.addr_out(config_seq_addr_out),
		.rd_data_out(config_data_out_shrt),
		.ren_out(config_seq_ren_out),
		.wen_out(config_seq_wen_out),
		.wr_data(config_seq_wr_data)
	);
endmodule
module LakeTop_W (
	clk,
	clk_en,
	config_addr_in,
	config_data_in,
	config_en,
	config_read,
	config_write,
	flush,
	input_width_16_num_0,
	input_width_16_num_1,
	input_width_16_num_2,
	input_width_16_num_3,
	input_width_1_num_0,
	input_width_1_num_1,
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality,
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0,
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1,
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2,
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3,
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4,
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5,
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable,
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr,
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0,
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1,
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2,
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3,
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4,
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_0,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_1,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_2,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_3,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_4,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_5,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_0,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_1,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_2,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_3,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_4,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_5,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_3,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_4,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_5,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_3,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_4,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_5,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_3,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_4,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_5,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_3,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_4,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_5,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_0,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_1,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_2,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_3,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_4,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_5,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_0,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_1,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_2,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_3,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_4,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_5,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4,
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4,
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5,
	mode,
	rst_n,
	tile_en,
	config_data_out,
	output_width_16_num_0,
	output_width_16_num_1,
	output_width_1_num_0,
	output_width_1_num_1,
	output_width_1_num_2
);
	input wire clk;
	input wire clk_en;
	input wire [7:0] config_addr_in;
	input wire [31:0] config_data_in;
	input wire config_en;
	input wire config_read;
	input wire config_write;
	input wire flush;
	input wire [15:0] input_width_16_num_0;
	input wire [15:0] input_width_16_num_1;
	input wire [15:0] input_width_16_num_2;
	input wire [15:0] input_width_16_num_3;
	input wire input_width_1_num_0;
	input wire input_width_1_num_1;
	input wire [3:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality;
	input wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0;
	input wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1;
	input wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2;
	input wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3;
	input wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4;
	input wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5;
	input wire mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable;
	input wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr;
	input wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0;
	input wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1;
	input wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2;
	input wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3;
	input wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4;
	input wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_0;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_1;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_2;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_3;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_4;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_5;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_0;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_1;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_2;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_3;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_4;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_5;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_3;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_4;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_5;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_3;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_4;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_5;
	input wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5;
	input wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_3;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_4;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_5;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_3;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_4;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_5;
	input wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5;
	input wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5;
	input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4;
	input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5;
	input wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_0;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_1;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_2;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_3;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_4;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_5;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_0;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_1;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_2;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_3;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_4;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_5;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4;
	input wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5;
	// input wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5;
	// input wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5;
	// input wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5;
	// input wire mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4;
	// input wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4;
	// input wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5;
	input wire [1:0] mode;
	input wire rst_n;
	input wire tile_en;
	output wire [31:0] config_data_out;
	output wire [15:0] output_width_16_num_0;
	output wire [15:0] output_width_16_num_1;
	output wire output_width_1_num_0;
	output wire output_width_1_num_1;
	output wire output_width_1_num_2;
	wire [95:0] LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges;
	wire [95:0] LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides;
	wire [23:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides;
	wire [23:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides;
	wire [23:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides;
	wire [23:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides;
	wire [95:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides;
	wire [95:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides;
	wire [95:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges;
	wire [95:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges;
	wire [95:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides;
	wire [95:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides;
	wire [95:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges;
	wire [95:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges;
	wire [47:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides;
	wire [47:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides;
	wire [47:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides;
	wire [47:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides;
	// wire [95:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges;
	// wire [95:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges;
	// wire [95:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides;
	// wire [95:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides;
	// wire [95:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges;
	// wire [95:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges;
	// wire [23:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides;
	// wire [23:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides;
	// wire [95:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides;
	// wire [95:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides;
	// wire [23:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides;
	// wire [23:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides;
	assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges[0+:16] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0;
	assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges[16+:16] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1;
	assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges[32+:16] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2;
	assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges[48+:16] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3;
	assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges[64+:16] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4;
	assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges[80+:16] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5;
	assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides[0+:16] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0;
	assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides[16+:16] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1;
	assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides[32+:16] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2;
	assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides[48+:16] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3;
	assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides[64+:16] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4;
	assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides[80+:16] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides[0+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_0;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides[4+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_1;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides[8+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_2;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides[12+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_3;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides[16+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_4;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides[20+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_5;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides[0+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_0;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides[4+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_1;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides[8+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_2;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides[12+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_3;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides[16+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_4;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides[20+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_5;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides[0+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides[4+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides[8+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides[12+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_3;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides[16+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_4;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides[20+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_5;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides[0+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides[4+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides[8+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides[12+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_3;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides[16+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_4;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides[20+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_5;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides[0+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides[16+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides[32+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides[48+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides[64+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides[80+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides[0+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides[16+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides[32+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides[48+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides[64+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides[80+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges[0+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges[16+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges[32+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges[48+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_3;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges[64+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_4;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges[80+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_5;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges[0+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges[16+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges[32+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges[48+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_3;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges[64+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_4;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges[80+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_5;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides[0+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides[16+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides[32+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides[48+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides[64+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides[80+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides[0+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides[16+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides[32+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides[48+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides[64+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides[80+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges[0+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges[16+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges[32+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges[48+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges[64+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges[80+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges[0+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges[16+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges[32+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges[48+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges[64+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges[80+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides[0+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_0;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides[8+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_1;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides[16+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_2;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides[24+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_3;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides[32+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_4;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides[40+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_5;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides[0+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_0;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides[8+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_1;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides[16+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_2;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides[24+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_3;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides[32+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_4;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides[40+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_5;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides[0+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides[8+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides[16+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides[24+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides[32+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides[40+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides[0+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides[8+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides[16+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides[24+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides[32+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4;
	assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides[40+:8] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges[0+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges[16+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges[32+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges[48+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges[64+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges[80+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges[0+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges[16+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges[32+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges[48+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges[64+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges[80+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides[0+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides[16+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides[32+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides[48+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides[64+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides[80+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides[0+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides[16+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides[32+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides[48+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides[64+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides[80+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges[0+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges[16+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges[32+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges[48+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges[64+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges[80+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges[0+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges[16+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges[32+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges[48+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges[64+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges[80+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides[0+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides[4+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides[8+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides[12+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides[16+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides[20+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides[0+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides[4+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides[8+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides[12+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides[16+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides[20+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides[0+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides[16+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides[32+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides[48+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides[64+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides[80+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides[0+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides[16+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides[32+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides[48+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides[64+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides[80+:16] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides[0+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides[4+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides[8+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides[12+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides[16+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides[20+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides[0+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides[4+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides[8+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides[12+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides[16+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4;
	// assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides[20+:4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5;
	LakeTop LakeTop(
		.clk(clk),
		.clk_en(clk_en),
		.config_addr_in(config_addr_in),
		.config_data_in(config_data_in),
		.config_en(config_en),
		.config_read(config_read),
		.config_write(config_write),
		.flush(flush),
		.input_width_16_num_0(input_width_16_num_0),
		.input_width_16_num_1(input_width_16_num_1),
		.input_width_16_num_2(input_width_16_num_2),
		.input_width_16_num_3(input_width_16_num_3),
		.input_width_1_num_0(input_width_1_num_0),
		.input_width_1_num_1(input_width_1_num_1),
		.mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality),
		.mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges(LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges),
		.mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable),
		.mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr),
		.mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides(LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides),
		.mode(mode),
		.rst_n(rst_n),
		.tile_en(tile_en),
		.config_data_out(config_data_out),
		.output_width_16_num_0(output_width_16_num_0),
		.output_width_16_num_1(output_width_16_num_1),
		.output_width_1_num_0(output_width_1_num_0),
		.output_width_1_num_1(output_width_1_num_1),
		.output_width_1_num_2(output_width_1_num_2)
	);
endmodule
module addr_gen_6_16 (
	clk,
	clk_en,
	flush,
	mux_sel,
	restart,
	rst_n,
	starting_addr,
	step,
	strides,
	addr_out
);
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire [2:0] mux_sel;
	input wire restart;
	input wire rst_n;
	input wire [15:0] starting_addr;
	input wire step;
	input wire [95:0] strides;
	output wire [15:0] addr_out;
	wire [15:0] calc_addr;
	reg [15:0] current_addr;
	wire [15:0] strt_addr;
	assign strt_addr = starting_addr;
	assign addr_out = calc_addr;
	assign calc_addr = strt_addr + current_addr;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			current_addr <= 16'h0000;
		else if (clk_en)
			if (flush)
				current_addr <= 16'h0000;
			else if (step)
				if (restart)
					current_addr <= 16'h0000;
				else
					current_addr <= current_addr + strides[mux_sel * 16+:16];
endmodule
module addr_gen_6_4 (
	clk,
	clk_en,
	flush,
	mux_sel,
	restart,
	rst_n,
	starting_addr,
	step,
	strides,
	addr_out
);
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire [2:0] mux_sel;
	input wire restart;
	input wire rst_n;
	input wire [3:0] starting_addr;
	input wire step;
	input wire [23:0] strides;
	output wire [3:0] addr_out;
	wire [3:0] calc_addr;
	reg [3:0] current_addr;
	wire [3:0] strt_addr;
	assign strt_addr = starting_addr;
	assign addr_out = calc_addr;
	assign calc_addr = strt_addr + current_addr;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			current_addr <= 4'h0;
		else if (clk_en)
			if (flush)
				current_addr <= 4'h0;
			else if (step)
				if (restart)
					current_addr <= 4'h0;
				else
					current_addr <= current_addr + strides[mux_sel * 4+:4];
endmodule
module addr_gen_6_8 (
	clk,
	clk_en,
	flush,
	mux_sel,
	restart,
	rst_n,
	starting_addr,
	step,
	strides,
	addr_out
);
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire [2:0] mux_sel;
	input wire restart;
	input wire rst_n;
	input wire [7:0] starting_addr;
	input wire step;
	input wire [47:0] strides;
	output wire [7:0] addr_out;
	wire [7:0] calc_addr;
	reg [7:0] current_addr;
	wire [7:0] strt_addr;
	assign strt_addr = starting_addr;
	assign addr_out = calc_addr;
	assign calc_addr = strt_addr + current_addr;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			current_addr <= 8'h00;
		else if (clk_en)
			if (flush)
				current_addr <= 8'h00;
			else if (step)
				if (restart)
					current_addr <= 8'h00;
				else
					current_addr <= current_addr + strides[mux_sel * 8+:8];
endmodule
module for_loop_6_16 (
	clk,
	clk_en,
	dimensionality,
	flush,
	ranges,
	rst_n,
	step,
	mux_sel_out,
	restart
);
	parameter CONFIG_WIDTH = 5'h10;
	parameter ITERATOR_SUPPORT = 4'h6;
	input wire clk;
	input wire clk_en;
	input wire [3:0] dimensionality;
	input wire flush;
	input wire [95:0] ranges;
	input wire rst_n;
	input wire step;
	output wire [2:0] mux_sel_out;
	output wire restart;
	reg [5:0] clear;
	reg [95:0] dim_counter;
	reg done;
	reg [5:0] inc;
	wire [15:0] inced_cnt;
	reg [5:0] max_value;
	wire maxed_value;
	reg [2:0] mux_sel;
	assign mux_sel_out = mux_sel;
	assign inced_cnt = dim_counter[mux_sel * 16+:16] + 16'h0001;
	assign maxed_value = (dim_counter[mux_sel * 16+:16] == ranges[mux_sel * 16+:16]) & inc[mux_sel];
	always @(*) begin
		mux_sel = 3'h0;
		done = 1'h0;
		if (~done)
			if (~max_value[0] & (dimensionality > 4'h0)) begin
				mux_sel = 3'h0;
				done = 1'h1;
			end
		if (~done)
			if (~max_value[1] & (dimensionality > 4'h1)) begin
				mux_sel = 3'h1;
				done = 1'h1;
			end
		if (~done)
			if (~max_value[2] & (dimensionality > 4'h2)) begin
				mux_sel = 3'h2;
				done = 1'h1;
			end
		if (~done)
			if (~max_value[3] & (dimensionality > 4'h3)) begin
				mux_sel = 3'h3;
				done = 1'h1;
			end
		if (~done)
			if (~max_value[4] & (dimensionality > 4'h4)) begin
				mux_sel = 3'h4;
				done = 1'h1;
			end
		if (~done)
			if (~max_value[5] & (dimensionality > 4'h5)) begin
				mux_sel = 3'h5;
				done = 1'h1;
			end
	end
	always @(*) begin
		clear[0] = 1'h0;
		if (((mux_sel > 3'h0) | ~done) & step)
			clear[0] = 1'h1;
	end
	always @(*) begin
		inc[0] = 1'h0;
		if (((5'h00 == 5'h00) & step) & (dimensionality > 4'h0))
			inc[0] = 1'h1;
		else if (((mux_sel == 3'h0) & step) & (dimensionality > 4'h0))
			inc[0] = 1'h1;
	end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			dim_counter[0+:16] <= 16'h0000;
		else if (clk_en)
			if (flush)
				dim_counter[0+:16] <= 16'h0000;
			else if (clear[0])
				dim_counter[0+:16] <= 16'h0000;
			else if (inc[0])
				dim_counter[0+:16] <= inced_cnt;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			max_value[0] <= 1'h0;
		else if (clk_en)
			if (flush)
				max_value[0] <= 1'h0;
			else if (clear[0])
				max_value[0] <= 1'h0;
			else if (inc[0])
				max_value[0] <= maxed_value;
	always @(*) begin
		clear[1] = 1'h0;
		if (((mux_sel > 3'h1) | ~done) & step)
			clear[1] = 1'h1;
	end
	always @(*) begin
		inc[1] = 1'h0;
		if (((5'h01 == 5'h00) & step) & (dimensionality > 4'h1))
			inc[1] = 1'h1;
		else if (((mux_sel == 3'h1) & step) & (dimensionality > 4'h1))
			inc[1] = 1'h1;
	end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			dim_counter[16+:16] <= 16'h0000;
		else if (clk_en)
			if (flush)
				dim_counter[16+:16] <= 16'h0000;
			else if (clear[1])
				dim_counter[16+:16] <= 16'h0000;
			else if (inc[1])
				dim_counter[16+:16] <= inced_cnt;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			max_value[1] <= 1'h0;
		else if (clk_en)
			if (flush)
				max_value[1] <= 1'h0;
			else if (clear[1])
				max_value[1] <= 1'h0;
			else if (inc[1])
				max_value[1] <= maxed_value;
	always @(*) begin
		clear[2] = 1'h0;
		if (((mux_sel > 3'h2) | ~done) & step)
			clear[2] = 1'h1;
	end
	always @(*) begin
		inc[2] = 1'h0;
		if (((5'h02 == 5'h00) & step) & (dimensionality > 4'h2))
			inc[2] = 1'h1;
		else if (((mux_sel == 3'h2) & step) & (dimensionality > 4'h2))
			inc[2] = 1'h1;
	end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			dim_counter[32+:16] <= 16'h0000;
		else if (clk_en)
			if (flush)
				dim_counter[32+:16] <= 16'h0000;
			else if (clear[2])
				dim_counter[32+:16] <= 16'h0000;
			else if (inc[2])
				dim_counter[32+:16] <= inced_cnt;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			max_value[2] <= 1'h0;
		else if (clk_en)
			if (flush)
				max_value[2] <= 1'h0;
			else if (clear[2])
				max_value[2] <= 1'h0;
			else if (inc[2])
				max_value[2] <= maxed_value;
	always @(*) begin
		clear[3] = 1'h0;
		if (((mux_sel > 3'h3) | ~done) & step)
			clear[3] = 1'h1;
	end
	always @(*) begin
		inc[3] = 1'h0;
		if (((5'h03 == 5'h00) & step) & (dimensionality > 4'h3))
			inc[3] = 1'h1;
		else if (((mux_sel == 3'h3) & step) & (dimensionality > 4'h3))
			inc[3] = 1'h1;
	end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			dim_counter[48+:16] <= 16'h0000;
		else if (clk_en)
			if (flush)
				dim_counter[48+:16] <= 16'h0000;
			else if (clear[3])
				dim_counter[48+:16] <= 16'h0000;
			else if (inc[3])
				dim_counter[48+:16] <= inced_cnt;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			max_value[3] <= 1'h0;
		else if (clk_en)
			if (flush)
				max_value[3] <= 1'h0;
			else if (clear[3])
				max_value[3] <= 1'h0;
			else if (inc[3])
				max_value[3] <= maxed_value;
	always @(*) begin
		clear[4] = 1'h0;
		if (((mux_sel > 3'h4) | ~done) & step)
			clear[4] = 1'h1;
	end
	always @(*) begin
		inc[4] = 1'h0;
		if (((5'h04 == 5'h00) & step) & (dimensionality > 4'h4))
			inc[4] = 1'h1;
		else if (((mux_sel == 3'h4) & step) & (dimensionality > 4'h4))
			inc[4] = 1'h1;
	end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			dim_counter[64+:16] <= 16'h0000;
		else if (clk_en)
			if (flush)
				dim_counter[64+:16] <= 16'h0000;
			else if (clear[4])
				dim_counter[64+:16] <= 16'h0000;
			else if (inc[4])
				dim_counter[64+:16] <= inced_cnt;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			max_value[4] <= 1'h0;
		else if (clk_en)
			if (flush)
				max_value[4] <= 1'h0;
			else if (clear[4])
				max_value[4] <= 1'h0;
			else if (inc[4])
				max_value[4] <= maxed_value;
	always @(*) begin
		clear[5] = 1'h0;
		if (((mux_sel > 3'h5) | ~done) & step)
			clear[5] = 1'h1;
	end
	always @(*) begin
		inc[5] = 1'h0;
		if (((5'h05 == 5'h00) & step) & (dimensionality > 4'h5))
			inc[5] = 1'h1;
		else if (((mux_sel == 3'h5) & step) & (dimensionality > 4'h5))
			inc[5] = 1'h1;
	end
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			dim_counter[80+:16] <= 16'h0000;
		else if (clk_en)
			if (flush)
				dim_counter[80+:16] <= 16'h0000;
			else if (clear[5])
				dim_counter[80+:16] <= 16'h0000;
			else if (inc[5])
				dim_counter[80+:16] <= inced_cnt;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			max_value[5] <= 1'h0;
		else if (clk_en)
			if (flush)
				max_value[5] <= 1'h0;
			else if (clear[5])
				max_value[5] <= 1'h0;
			else if (inc[5])
				max_value[5] <= maxed_value;
	assign restart = step & ~done;
endmodule
module sched_gen_6_16 (
	clk,
	clk_en,
	cycle_count,
	enable,
	finished,
	flush,
	mux_sel,
	rst_n,
	sched_addr_gen_starting_addr,
	sched_addr_gen_strides,
	valid_output
);
	input wire clk;
	input wire clk_en;
	input wire [15:0] cycle_count;
	input wire enable;
	input wire finished;
	input wire flush;
	input wire [2:0] mux_sel;
	input wire rst_n;
	input wire [15:0] sched_addr_gen_starting_addr;
	input wire [95:0] sched_addr_gen_strides;
	output reg valid_output;
	wire [15:0] addr_out;
	wire valid_gate;
	reg valid_gate_inv;
	reg valid_out;
	assign valid_gate = ~valid_gate_inv;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			valid_gate_inv <= 1'h0;
		else if (clk_en)
			if (flush)
				valid_gate_inv <= 1'h0;
			else if (finished)
				valid_gate_inv <= 1'h1;
	always @(*) valid_out = ((cycle_count == addr_out) & valid_gate) & enable;
	always @(*) valid_output = valid_out;
	addr_gen_6_16 sched_addr_gen(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(mux_sel),
		.restart(1'h0),
		.rst_n(rst_n),
		.starting_addr(sched_addr_gen_starting_addr),
		.step(valid_out),
		.strides(sched_addr_gen_strides),
		.addr_out(addr_out)
	);
endmodule
module sram_idk_0 (
	clk,
	clk_en,
	data_in_p0,
	flush,
	read_addr_p0,
	read_addr_p1,
	read_enable_p0,
	read_enable_p1,
	write_addr_p0,
	write_enable_p0,
	data_out_p0,
	data_out_p1
);
	input wire clk;
	input wire clk_en;
	input wire [31:0] data_in_p0;
	input wire flush;
	input wire [7:0] read_addr_p0;
	input wire [7:0] read_addr_p1;
	input wire read_enable_p0;
	input wire read_enable_p1;
	input wire [7:0] write_addr_p0;
	input wire write_enable_p0;
	output reg [31:0] data_out_p0;
	output reg [31:0] data_out_p1;
	reg [31:0] data_array [255:0];
	always @(posedge clk)
		if (clk_en)
			if (write_enable_p0 == 1'h1)
				data_array[write_addr_p0] <= data_in_p0;
			else if (read_enable_p0)
				data_out_p0 <= data_array[read_addr_p0];
	always @(posedge clk)
		if (clk_en)
			if (read_enable_p1 == 1'h1)
				data_out_p1 <= data_array[read_addr_p1];
endmodule
module stencil_valid (
	clk,
	clk_en,
	flush,
	loops_stencil_valid_dimensionality,
	loops_stencil_valid_ranges,
	rst_n,
	stencil_valid_sched_gen_enable,
	stencil_valid_sched_gen_sched_addr_gen_starting_addr,
	stencil_valid_sched_gen_sched_addr_gen_strides,
	stencil_valid
);
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire [3:0] loops_stencil_valid_dimensionality;
	input wire [95:0] loops_stencil_valid_ranges;
	input wire rst_n;
	input wire stencil_valid_sched_gen_enable;
	input wire [15:0] stencil_valid_sched_gen_sched_addr_gen_starting_addr;
	input wire [95:0] stencil_valid_sched_gen_sched_addr_gen_strides;
	output wire stencil_valid;
	reg [15:0] cycle_count;
	wire [2:0] loops_stencil_valid_mux_sel_out;
	wire loops_stencil_valid_restart;
	wire stencil_valid_internal;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			cycle_count <= 16'h0000;
		else if (clk_en)
			if (flush)
				cycle_count <= 16'h0000;
			else
				cycle_count <= cycle_count + 16'h0001;
	assign stencil_valid = stencil_valid_internal;
	for_loop_6_16 #(
		.CONFIG_WIDTH(5'h10),
		.ITERATOR_SUPPORT(4'h6)
	) loops_stencil_valid(
		.clk(clk),
		.clk_en(clk_en),
		.dimensionality(loops_stencil_valid_dimensionality),
		.flush(flush),
		.ranges(loops_stencil_valid_ranges),
		.rst_n(rst_n),
		.step(stencil_valid_internal),
		.mux_sel_out(loops_stencil_valid_mux_sel_out),
		.restart(loops_stencil_valid_restart)
	);
	sched_gen_6_16 stencil_valid_sched_gen(
		.clk(clk),
		.clk_en(clk_en),
		.cycle_count(cycle_count),
		.enable(stencil_valid_sched_gen_enable),
		.finished(loops_stencil_valid_restart),
		.flush(flush),
		.mux_sel(loops_stencil_valid_mux_sel_out),
		.rst_n(rst_n),
		.sched_addr_gen_starting_addr(stencil_valid_sched_gen_sched_addr_gen_starting_addr),
		.sched_addr_gen_strides(stencil_valid_sched_gen_sched_addr_gen_strides),
		.valid_output(stencil_valid_internal)
	);
endmodule
module stencil_valid_flat (
	clk,
	clk_en,
	flush,
	rst_n,
	stencil_valid_inst_loops_stencil_valid_dimensionality,
	stencil_valid_inst_loops_stencil_valid_ranges,
	stencil_valid_inst_stencil_valid_sched_gen_enable,
	stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr,
	stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides,
	stencil_valid_f_
);
	input wire clk;
	input wire clk_en;
	input wire flush;
	input wire rst_n;
	input wire [3:0] stencil_valid_inst_loops_stencil_valid_dimensionality;
	input wire [95:0] stencil_valid_inst_loops_stencil_valid_ranges;
	input wire stencil_valid_inst_stencil_valid_sched_gen_enable;
	input wire [15:0] stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr;
	input wire [95:0] stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides;
	output wire stencil_valid_f_;
	stencil_valid stencil_valid_inst(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.loops_stencil_valid_dimensionality(stencil_valid_inst_loops_stencil_valid_dimensionality),
		.loops_stencil_valid_ranges(stencil_valid_inst_loops_stencil_valid_ranges),
		.rst_n(rst_n),
		.stencil_valid_sched_gen_enable(stencil_valid_inst_stencil_valid_sched_gen_enable),
		.stencil_valid_sched_gen_sched_addr_gen_starting_addr(stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr),
		.stencil_valid_sched_gen_sched_addr_gen_strides(stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides),
		.stencil_valid(stencil_valid_f_)
	);
endmodule
module storage_config_seq (
	clk,
	clk_en,
	config_addr_in,
	config_data_in,
	config_en,
	config_rd,
	config_wr,
	flush,
	rd_data_stg,
	rst_n,
	addr_out,
	rd_data_out,
	ren_out,
	wen_out,
	wr_data
);
	input wire clk;
	input wire clk_en;
	input wire [7:0] config_addr_in;
	input wire [15:0] config_data_in;
	input wire config_en;
	input wire config_rd;
	input wire config_wr;
	input wire flush;
	input wire [31:0] rd_data_stg;
	input wire rst_n;
	output wire [7:0] addr_out;
	output wire [15:0] rd_data_out;
	output wire ren_out;
	output wire wen_out;
	output wire [31:0] wr_data;
	reg cnt;
	reg [15:0] data_wr_reg;
	reg rd_cnt;
	assign addr_out = config_addr_in[7:0];
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			cnt <= 1'h0;
		else if (flush)
			cnt <= 1'h0;
		else if ((config_wr | config_rd) & |config_en)
			cnt <= cnt + 1'h1;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			rd_cnt <= 1'h0;
		else if (flush)
			rd_cnt <= 1'h0;
		else
			rd_cnt <= cnt;
	assign rd_data_out[0+:16] = rd_data_stg[rd_cnt * 16+:16];
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			data_wr_reg <= 16'h0000;
		else if (flush)
			data_wr_reg <= 16'h0000;
		else if (config_wr & (cnt < 1'h1))
			data_wr_reg[cnt * 16+:16] <= config_data_in;
	assign wr_data[0+:16] = data_wr_reg[0+:16];
	assign wr_data[16+:16] = config_data_in;
	assign wen_out = config_wr & (cnt == 1'h1);
	assign ren_out = config_rd;
endmodule
module strg_ram (
	clk,
	clk_en,
	data_from_strg,
	data_in,
	flush,
	rd_addr_in,
	ren,
	rst_n,
	wen,
	wr_addr_in,
	addr_out,
	data_out,
	data_to_strg,
	ready,
	ren_to_strg,
	valid_out,
	wen_to_strg
);
	input wire clk;
	input wire clk_en;
	input wire [31:0] data_from_strg;
	input wire [15:0] data_in;
	input wire flush;
	input wire [15:0] rd_addr_in;
	input wire ren;
	input wire rst_n;
	input wire wen;
	input wire [15:0] wr_addr_in;
	output reg [7:0] addr_out;
	output reg [15:0] data_out;
	output wire [31:0] data_to_strg;
	output reg ready;
	output wire ren_to_strg;
	output reg valid_out;
	output wire wen_to_strg;
	reg [15:0] addr_to_write;
	reg [31:0] data_combined;
	reg [15:0] data_to_write;
	reg [1:0] r_w_seq_current_state;
	reg [1:0] r_w_seq_next_state;
	wire [15:0] rd_addr;
	wire rd_bank;
	reg read_gate;
	wire [15:0] wr_addr;
	reg write_gate;
	assign wr_addr = wr_addr_in;
	assign rd_addr = rd_addr_in;
	assign rd_bank = 1'h0;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			data_to_write <= 16'h0000;
		else if (clk_en)
			if (flush)
				data_to_write <= 16'h0000;
			else
				data_to_write <= data_in;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			addr_to_write <= 16'h0000;
		else if (clk_en)
			if (flush)
				addr_to_write <= 16'h0000;
			else
				addr_to_write <= wr_addr;
	assign data_to_strg[0+:32] = data_combined;
	assign ren_to_strg = (wen | ren) & read_gate;
	assign wen_to_strg = write_gate;
	always @(*) begin
		addr_out[0+:8] = rd_addr[8:1];
		if (wen & ~write_gate)
			addr_out[0+:8] = wr_addr[8:1];
		else if (write_gate)
			addr_out[0+:8] = addr_to_write[8:1];
	end
	always @(*)
		if (addr_to_write[0] == 1'h0)
			data_combined[0+:16] = data_to_write;
		else
			data_combined[0+:16] = data_from_strg[(rd_bank * 2) * 16+:16];
	always @(*)
		if (addr_to_write[0] == 1'h1)
			data_combined[16+:16] = data_to_write;
		else
			data_combined[16+:16] = data_from_strg[((rd_bank * 2) + 1) * 16+:16];
	localparam [1:0] IDLE = 2'h0;
	always @(posedge clk or negedge rst_n)
		if (!rst_n)
			r_w_seq_current_state <= IDLE;
		else
			r_w_seq_current_state <= r_w_seq_next_state;
	localparam [1:0] MODIFY = 2'h1;
	localparam [1:0] READ = 2'h2;
	localparam [1:0] _DEFAULT = 2'h3;
	always @(*) begin
		r_w_seq_next_state = r_w_seq_current_state;
		case (r_w_seq_current_state)
			IDLE:
				if (~wen & ~ren)
					r_w_seq_next_state = IDLE;
				else if (wen)
					r_w_seq_next_state = MODIFY;
				else if (ren & ~wen)
					r_w_seq_next_state = READ;
			MODIFY: r_w_seq_next_state = IDLE;
			READ:
				if (~wen & ~ren)
					r_w_seq_next_state = IDLE;
				else if (wen)
					r_w_seq_next_state = MODIFY;
				else if (ren & ~wen)
					r_w_seq_next_state = READ;
			_DEFAULT: r_w_seq_next_state = _DEFAULT;
		endcase
	end
	always @(*)
		case (r_w_seq_current_state)
			IDLE: begin : r_w_seq_IDLE_Output
				data_out = 16'h0000;
				read_gate = 1'h1;
				ready = 1'h1;
				valid_out = 1'h0;
				write_gate = 1'h0;
			end
			MODIFY: begin : r_w_seq_MODIFY_Output
				data_out = 16'h0000;
				read_gate = 1'h0;
				ready = 1'h0;
				valid_out = 1'h0;
				write_gate = 1'h1;
			end
			READ: begin : r_w_seq_READ_Output
				data_out = data_from_strg[((rd_bank * 2) + addr_to_write[0]) * 16+:16];
				read_gate = 1'h1;
				ready = 1'h1;
				valid_out = 1'h1;
				write_gate = 1'h0;
			end
			_DEFAULT: begin : r_w_seq__DEFAULT_Output
				data_out = 16'h0000;
				read_gate = 1'h0;
				ready = 1'h0;
				valid_out = 1'h0;
				write_gate = 1'h0;
			end
		endcase
endmodule
module strg_ram_flat (
	clk,
	clk_en,
	data_from_strg_lifted,
	data_in_f_,
	flush,
	rd_addr_in_f_,
	ren_f_,
	rst_n,
	wen_f_,
	wr_addr_in_f_,
	addr_out_lifted,
	data_out_f_,
	data_to_strg_lifted,
	ready_f_,
	ren_to_strg_lifted,
	valid_out_f_,
	wen_to_strg_lifted
);
	input wire clk;
	input wire clk_en;
	input wire [31:0] data_from_strg_lifted;
	input wire [15:0] data_in_f_;
	input wire flush;
	input wire [15:0] rd_addr_in_f_;
	input wire ren_f_;
	input wire rst_n;
	input wire wen_f_;
	input wire [15:0] wr_addr_in_f_;
	output wire [7:0] addr_out_lifted;
	output wire [15:0] data_out_f_;
	output wire [31:0] data_to_strg_lifted;
	output wire ready_f_;
	output wire ren_to_strg_lifted;
	output wire valid_out_f_;
	output wire wen_to_strg_lifted;
	wire [15:0] data_in_f__intercept;
	wire [15:0] data_out_f__intercept;
	wire [15:0] rd_addr_in_f__intercept;
	wire [15:0] strg_ram_inst_data_in;
	wire [15:0] strg_ram_inst_data_out;
	wire [15:0] strg_ram_inst_rd_addr_in;
	wire [15:0] strg_ram_inst_wr_addr_in;
	wire [15:0] wr_addr_in_f__intercept;
	assign strg_ram_inst_rd_addr_in = rd_addr_in_f__intercept[0+:16];
	assign rd_addr_in_f__intercept = rd_addr_in_f_;
	assign strg_ram_inst_data_in = data_in_f__intercept[0+:16];
	assign data_in_f__intercept = data_in_f_;
	assign strg_ram_inst_wr_addr_in = wr_addr_in_f__intercept[0+:16];
	assign wr_addr_in_f__intercept = wr_addr_in_f_;
	assign data_out_f__intercept[0+:16] = strg_ram_inst_data_out;
	assign data_out_f_ = data_out_f__intercept;
	strg_ram strg_ram_inst(
		.clk(clk),
		.clk_en(clk_en),
		.data_from_strg(data_from_strg_lifted),
		.data_in(strg_ram_inst_data_in),
		.flush(flush),
		.rd_addr_in(strg_ram_inst_rd_addr_in),
		.ren(ren_f_),
		.rst_n(rst_n),
		.wen(wen_f_),
		.wr_addr_in(strg_ram_inst_wr_addr_in),
		.addr_out(addr_out_lifted),
		.data_out(strg_ram_inst_data_out),
		.data_to_strg(data_to_strg_lifted),
		.ready(ready_f_),
		.ren_to_strg(ren_to_strg_lifted),
		.valid_out(valid_out_f_),
		.wen_to_strg(wen_to_strg_lifted)
	);
endmodule
module strg_ub_agg_only (
	agg_read,
	agg_read_addr_gen_0_starting_addr,
	agg_read_addr_gen_0_strides,
	agg_read_addr_gen_1_starting_addr,
	agg_read_addr_gen_1_strides,
	agg_write_addr_gen_0_starting_addr,
	agg_write_addr_gen_0_strides,
	agg_write_addr_gen_1_starting_addr,
	agg_write_addr_gen_1_strides,
	agg_write_sched_gen_0_enable,
	agg_write_sched_gen_0_sched_addr_gen_starting_addr,
	agg_write_sched_gen_0_sched_addr_gen_strides,
	agg_write_sched_gen_1_enable,
	agg_write_sched_gen_1_sched_addr_gen_starting_addr,
	agg_write_sched_gen_1_sched_addr_gen_strides,
	clk,
	clk_en,
	cycle_count,
	data_in,
	floop_mux_sel,
	floop_restart,
	flush,
	loops_in2buf_0_dimensionality,
	loops_in2buf_0_ranges,
	loops_in2buf_1_dimensionality,
	loops_in2buf_1_ranges,
	rst_n,
	agg_data_out
);
	input wire [1:0] agg_read;
	input wire [3:0] agg_read_addr_gen_0_starting_addr;
	input wire [23:0] agg_read_addr_gen_0_strides;
	input wire [3:0] agg_read_addr_gen_1_starting_addr;
	input wire [23:0] agg_read_addr_gen_1_strides;
	input wire [3:0] agg_write_addr_gen_0_starting_addr;
	input wire [23:0] agg_write_addr_gen_0_strides;
	input wire [3:0] agg_write_addr_gen_1_starting_addr;
	input wire [23:0] agg_write_addr_gen_1_strides;
	input wire agg_write_sched_gen_0_enable;
	input wire [15:0] agg_write_sched_gen_0_sched_addr_gen_starting_addr;
	input wire [95:0] agg_write_sched_gen_0_sched_addr_gen_strides;
	input wire agg_write_sched_gen_1_enable;
	input wire [15:0] agg_write_sched_gen_1_sched_addr_gen_starting_addr;
	input wire [95:0] agg_write_sched_gen_1_sched_addr_gen_strides;
	input wire clk;
	input wire clk_en;
	input wire [15:0] cycle_count;
	input wire [31:0] data_in;
	input wire [5:0] floop_mux_sel;
	input wire [1:0] floop_restart;
	input wire flush;
	input wire [3:0] loops_in2buf_0_dimensionality;
	input wire [95:0] loops_in2buf_0_ranges;
	input wire [3:0] loops_in2buf_1_dimensionality;
	input wire [95:0] loops_in2buf_1_ranges;
	input wire rst_n;
	output reg [63:0] agg_data_out;
	// reg [255:0] agg;
	reg [255:0] agg0;  // 通道0使用的寄存器 
	reg [255:0] agg1;  // 通道1使用的寄存器
	wire [3:0] agg_read_addr;
	wire [3:0] agg_read_addr_gen_0_addr_out;
	wire [2:0] agg_read_addr_gen_0_mux_sel;
	wire agg_read_addr_gen_0_restart;
	wire agg_read_addr_gen_0_step;
	wire [3:0] agg_read_addr_gen_1_addr_out;
	wire [2:0] agg_read_addr_gen_1_mux_sel;
	wire agg_read_addr_gen_1_restart;
	wire agg_read_addr_gen_1_step;
	wire [15:0] agg_read_addr_gen_out;
	wire [1:0] agg_write;
	wire [5:0] agg_write_addr;
	wire [3:0] agg_write_addr_gen_0_addr_out;
	wire agg_write_addr_gen_0_step;
	wire [3:0] agg_write_addr_gen_1_addr_out;
	wire agg_write_addr_gen_1_step;
	wire agg_write_sched_gen_0_valid_output;
	wire agg_write_sched_gen_1_valid_output;
	wire [2:0] loops_in2buf_0_mux_sel_out;
	wire loops_in2buf_0_restart;
	wire loops_in2buf_0_step;
	wire [2:0] loops_in2buf_1_mux_sel_out;
	wire loops_in2buf_1_restart;
	wire loops_in2buf_1_step;
	assign loops_in2buf_0_step = agg_write[0];
	assign agg_write_addr_gen_0_step = agg_write[0];
	assign agg_write_addr[0+:3] = agg_write_addr_gen_0_addr_out[2:0];
	assign agg_write[0] = agg_write_sched_gen_0_valid_output;
	// always @(posedge clk)
	// 	if (clk_en)
	// 		if (agg_write[0])
	// 			agg[((agg_write_addr[2-:2] * 2) + agg_write_addr[0]) * 16+:16] <= data_in[0+:16];
	assign agg_read_addr_gen_0_step = agg_read[0];
	assign agg_read_addr_gen_0_restart = floop_restart[0];
	assign agg_read_addr_gen_0_mux_sel = floop_mux_sel[0+:3];
	assign agg_read_addr_gen_out[3-:4] = agg_read_addr_gen_0_addr_out;
	assign agg_read_addr_gen_out[7-:4] = 4'h0;
	assign agg_read_addr[0+:2] = agg_read_addr_gen_out[1-:2];
	// always @(*) agg_data_out[0+:32] = agg[16 * (agg_read_addr[0+:2] * 2)+:32];
	assign loops_in2buf_1_step = agg_write[1];
	assign agg_write_addr_gen_1_step = agg_write[1];
	assign agg_write_addr[3+:3] = agg_write_addr_gen_1_addr_out[2:0];
	assign agg_write[1] = agg_write_sched_gen_1_valid_output;
	// always @(posedge clk)
	// 	if (clk_en)
	// 		if (agg_write[1])
	// 			agg[(((4 + agg_write_addr[5-:2]) * 2) + agg_write_addr[3]) * 16+:16] <= data_in[16+:16];
	assign agg_read_addr_gen_1_step = agg_read[1];
	assign agg_read_addr_gen_1_restart = floop_restart[1];
	assign agg_read_addr_gen_1_mux_sel = floop_mux_sel[3+:3];
	assign agg_read_addr_gen_out[11-:4] = agg_read_addr_gen_1_addr_out;
	assign agg_read_addr_gen_out[15-:4] = 4'h0;
	assign agg_read_addr[2+:2] = agg_read_addr_gen_out[9-:2];
	// always @(*) agg_data_out[32+:32] = agg[16 * ((4 + agg_read_addr[2+:2]) * 2)+:32];
	
	// 通道0写入agg0
	always @(posedge clk) begin
		if (!rst_n) begin
			agg0 <= 256'b0;
		end
		else if (clk_en && agg_write[0]) begin
			agg0[((agg_write_addr[2-:2] * 2) + agg_write_addr[0]) * 16+:16] <= data_in[0+:16];
		end
	end

	// 通道1写入agg1
	always @(posedge clk) begin
		if (!rst_n) begin
			agg1 <= 256'b0;
		end
		else if (clk_en && agg_write[1]) begin
			agg1[(((4 + agg_write_addr[5-:2]) * 2) + agg_write_addr[3]) * 16+:16] <= data_in[16+:16];
		end
	end

	// 读取逻辑也需要修改
	always @(*) begin
		agg_data_out[0+:32] = agg0[16 * (agg_read_addr[0+:2] * 2)+:32];
		agg_data_out[32+:32] = agg1[16 * ((4 + agg_read_addr[2+:2]) * 2)+:32];
	end
	
	for_loop_6_16 #(
		.CONFIG_WIDTH(5'h10),
		.ITERATOR_SUPPORT(4'h6)
	) loops_in2buf_0(
		.clk(clk),
		.clk_en(clk_en),
		.dimensionality(loops_in2buf_0_dimensionality),
		.flush(flush),
		.ranges(loops_in2buf_0_ranges),
		.rst_n(rst_n),
		.step(loops_in2buf_0_step),
		.mux_sel_out(loops_in2buf_0_mux_sel_out),
		.restart(loops_in2buf_0_restart)
	);
	addr_gen_6_4 agg_write_addr_gen_0(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(loops_in2buf_0_mux_sel_out),
		.restart(loops_in2buf_0_restart),
		.rst_n(rst_n),
		.starting_addr(agg_write_addr_gen_0_starting_addr),
		.step(agg_write_addr_gen_0_step),
		.strides(agg_write_addr_gen_0_strides),
		.addr_out(agg_write_addr_gen_0_addr_out)
	);
	sched_gen_6_16 agg_write_sched_gen_0(
		.clk(clk),
		.clk_en(clk_en),
		.cycle_count(cycle_count),
		.enable(agg_write_sched_gen_0_enable),
		.finished(loops_in2buf_0_restart),
		.flush(flush),
		.mux_sel(loops_in2buf_0_mux_sel_out),
		.rst_n(rst_n),
		.sched_addr_gen_starting_addr(agg_write_sched_gen_0_sched_addr_gen_starting_addr),
		.sched_addr_gen_strides(agg_write_sched_gen_0_sched_addr_gen_strides),
		.valid_output(agg_write_sched_gen_0_valid_output)
	);
	addr_gen_6_4 agg_read_addr_gen_0(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(agg_read_addr_gen_0_mux_sel),
		.restart(agg_read_addr_gen_0_restart),
		.rst_n(rst_n),
		.starting_addr(agg_read_addr_gen_0_starting_addr),
		.step(agg_read_addr_gen_0_step),
		.strides(agg_read_addr_gen_0_strides),
		.addr_out(agg_read_addr_gen_0_addr_out)
	);
	for_loop_6_16 #(
		.CONFIG_WIDTH(5'h10),
		.ITERATOR_SUPPORT(4'h6)
	) loops_in2buf_1(
		.clk(clk),
		.clk_en(clk_en),
		.dimensionality(loops_in2buf_1_dimensionality),
		.flush(flush),
		.ranges(loops_in2buf_1_ranges),
		.rst_n(rst_n),
		.step(loops_in2buf_1_step),
		.mux_sel_out(loops_in2buf_1_mux_sel_out),
		.restart(loops_in2buf_1_restart)
	);
	addr_gen_6_4 agg_write_addr_gen_1(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(loops_in2buf_1_mux_sel_out),
		.restart(loops_in2buf_1_restart),
		.rst_n(rst_n),
		.starting_addr(agg_write_addr_gen_1_starting_addr),
		.step(agg_write_addr_gen_1_step),
		.strides(agg_write_addr_gen_1_strides),
		.addr_out(agg_write_addr_gen_1_addr_out)
	);
	sched_gen_6_16 agg_write_sched_gen_1(
		.clk(clk),
		.clk_en(clk_en),
		.cycle_count(cycle_count),
		.enable(agg_write_sched_gen_1_enable),
		.finished(loops_in2buf_1_restart),
		.flush(flush),
		.mux_sel(loops_in2buf_1_mux_sel_out),
		.rst_n(rst_n),
		.sched_addr_gen_starting_addr(agg_write_sched_gen_1_sched_addr_gen_starting_addr),
		.sched_addr_gen_strides(agg_write_sched_gen_1_sched_addr_gen_strides),
		.valid_output(agg_write_sched_gen_1_valid_output)
	);
	addr_gen_6_4 agg_read_addr_gen_1(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(agg_read_addr_gen_1_mux_sel),
		.restart(agg_read_addr_gen_1_restart),
		.rst_n(rst_n),
		.starting_addr(agg_read_addr_gen_1_starting_addr),
		.step(agg_read_addr_gen_1_step),
		.strides(agg_read_addr_gen_1_strides),
		.addr_out(agg_read_addr_gen_1_addr_out)
	);
endmodule
module strg_ub_agg_sram_shared (
	agg_read_sched_gen_0_enable,
	agg_read_sched_gen_0_sched_addr_gen_starting_addr,
	agg_read_sched_gen_0_sched_addr_gen_strides,
	agg_read_sched_gen_1_enable,
	agg_read_sched_gen_1_sched_addr_gen_starting_addr,
	agg_read_sched_gen_1_sched_addr_gen_strides,
	clk,
	clk_en,
	cycle_count,
	flush,
	loops_in2buf_autovec_write_0_dimensionality,
	loops_in2buf_autovec_write_0_ranges,
	loops_in2buf_autovec_write_1_dimensionality,
	loops_in2buf_autovec_write_1_ranges,
	rst_n,
	agg_read_out,
	floop_mux_sel,
	floop_restart
);
	input wire agg_read_sched_gen_0_enable;
	input wire [15:0] agg_read_sched_gen_0_sched_addr_gen_starting_addr;
	input wire [95:0] agg_read_sched_gen_0_sched_addr_gen_strides;
	input wire agg_read_sched_gen_1_enable;
	input wire [15:0] agg_read_sched_gen_1_sched_addr_gen_starting_addr;
	input wire [95:0] agg_read_sched_gen_1_sched_addr_gen_strides;
	input wire clk;
	input wire clk_en;
	input wire [15:0] cycle_count;
	input wire flush;
	input wire [3:0] loops_in2buf_autovec_write_0_dimensionality;
	input wire [95:0] loops_in2buf_autovec_write_0_ranges;
	input wire [3:0] loops_in2buf_autovec_write_1_dimensionality;
	input wire [95:0] loops_in2buf_autovec_write_1_ranges;
	input wire rst_n;
	output wire [1:0] agg_read_out;
	output wire [5:0] floop_mux_sel;
	output wire [1:0] floop_restart;
	wire [1:0] agg_read;
	wire agg_read_sched_gen_0_valid_output;
	wire agg_read_sched_gen_1_valid_output;
	wire [2:0] loops_in2buf_autovec_write_0_mux_sel_out;
	wire loops_in2buf_autovec_write_0_restart;
	wire loops_in2buf_autovec_write_0_step;
	wire [2:0] loops_in2buf_autovec_write_1_mux_sel_out;
	wire loops_in2buf_autovec_write_1_restart;
	wire loops_in2buf_autovec_write_1_step;
	assign agg_read_out = agg_read;
	assign loops_in2buf_autovec_write_0_step = agg_read[0];
	assign floop_mux_sel[0+:3] = loops_in2buf_autovec_write_0_mux_sel_out;
	assign floop_restart[0] = loops_in2buf_autovec_write_0_restart;
	assign agg_read[0] = agg_read_sched_gen_0_valid_output;
	assign loops_in2buf_autovec_write_1_step = agg_read[1];
	assign floop_mux_sel[3+:3] = loops_in2buf_autovec_write_1_mux_sel_out;
	assign floop_restart[1] = loops_in2buf_autovec_write_1_restart;
	assign agg_read[1] = agg_read_sched_gen_1_valid_output;
	for_loop_6_16 #(
		.CONFIG_WIDTH(5'h10),
		.ITERATOR_SUPPORT(4'h6)
	) loops_in2buf_autovec_write_0(
		.clk(clk),
		.clk_en(clk_en),
		.dimensionality(loops_in2buf_autovec_write_0_dimensionality),
		.flush(flush),
		.ranges(loops_in2buf_autovec_write_0_ranges),
		.rst_n(rst_n),
		.step(loops_in2buf_autovec_write_0_step),
		.mux_sel_out(loops_in2buf_autovec_write_0_mux_sel_out),
		.restart(loops_in2buf_autovec_write_0_restart)
	);
	sched_gen_6_16 agg_read_sched_gen_0(
		.clk(clk),
		.clk_en(clk_en),
		.cycle_count(cycle_count),
		.enable(agg_read_sched_gen_0_enable),
		.finished(loops_in2buf_autovec_write_0_restart),
		.flush(flush),
		.mux_sel(loops_in2buf_autovec_write_0_mux_sel_out),
		.rst_n(rst_n),
		.sched_addr_gen_starting_addr(agg_read_sched_gen_0_sched_addr_gen_starting_addr),
		.sched_addr_gen_strides(agg_read_sched_gen_0_sched_addr_gen_strides),
		.valid_output(agg_read_sched_gen_0_valid_output)
	);
	for_loop_6_16 #(
		.CONFIG_WIDTH(5'h10),
		.ITERATOR_SUPPORT(4'h6)
	) loops_in2buf_autovec_write_1(
		.clk(clk),
		.clk_en(clk_en),
		.dimensionality(loops_in2buf_autovec_write_1_dimensionality),
		.flush(flush),
		.ranges(loops_in2buf_autovec_write_1_ranges),
		.rst_n(rst_n),
		.step(loops_in2buf_autovec_write_1_step),
		.mux_sel_out(loops_in2buf_autovec_write_1_mux_sel_out),
		.restart(loops_in2buf_autovec_write_1_restart)
	);
	sched_gen_6_16 agg_read_sched_gen_1(
		.clk(clk),
		.clk_en(clk_en),
		.cycle_count(cycle_count),
		.enable(agg_read_sched_gen_1_enable),
		.finished(loops_in2buf_autovec_write_1_restart),
		.flush(flush),
		.mux_sel(loops_in2buf_autovec_write_1_mux_sel_out),
		.rst_n(rst_n),
		.sched_addr_gen_starting_addr(agg_read_sched_gen_1_sched_addr_gen_starting_addr),
		.sched_addr_gen_strides(agg_read_sched_gen_1_sched_addr_gen_strides),
		.valid_output(agg_read_sched_gen_1_valid_output)
	);
endmodule
module strg_ub_sram_only (
	agg_data_out,
	agg_read,
	clk,
	clk_en,
	cycle_count,
	floop_mux_sel,
	floop_restart,
	flush,
	input_addr_gen_0_starting_addr,
	input_addr_gen_0_strides,
	input_addr_gen_1_starting_addr,
	input_addr_gen_1_strides,
	// loops_sram2tb_mux_sel,
	// loops_sram2tb_restart,
	output_addr_gen_0_starting_addr,
	output_addr_gen_0_strides,
	output_addr_gen_1_starting_addr,
	output_addr_gen_1_strides,
	rst_n,
	t_read,
	data_to_sram,
	rd_addr_to_sram,
	ren_to_sram,
	wen_to_sram,
	wr_addr_to_sram
);
	input wire [63:0] agg_data_out;
	input wire [1:0] agg_read;
	input wire clk;
	input wire clk_en;
	input wire [15:0] cycle_count;
	input wire [5:0] floop_mux_sel;
	input wire [1:0] floop_restart;
	input wire flush;
	input wire [7:0] input_addr_gen_0_starting_addr;
	input wire [47:0] input_addr_gen_0_strides;
	input wire [7:0] input_addr_gen_1_starting_addr;
	input wire [47:0] input_addr_gen_1_strides;
	// input wire [5:0] loops_sram2tb_mux_sel;
	// input wire [1:0] loops_sram2tb_restart;
	input wire [7:0] output_addr_gen_0_starting_addr;
	input wire [47:0] output_addr_gen_0_strides;
	input wire [7:0] output_addr_gen_1_starting_addr;
	input wire [47:0] output_addr_gen_1_strides;
	input wire rst_n;
	input wire [1:0] t_read;
	output wire [31:0] data_to_sram;
	output wire [7:0] rd_addr_to_sram;
	output wire ren_to_sram;
	output wire wen_to_sram;
	output wire [7:0] wr_addr_to_sram;
	reg [31:0] decode_ret_agg_read_agg_data_out;
	reg [15:0] decode_ret_agg_read_s_write_addr;
	reg [15:0] decode_ret_t_read_s_read_addr;
	reg decode_sel_done_agg_read_agg_data_out;
	reg decode_sel_done_agg_read_s_write_addr;
	reg decode_sel_done_t_read_s_read_addr;
	wire [7:0] input_addr_gen_0_addr_out;
	wire [2:0] input_addr_gen_0_mux_sel;
	wire input_addr_gen_0_restart;
	wire input_addr_gen_0_step;
	wire [7:0] input_addr_gen_1_addr_out;
	wire [2:0] input_addr_gen_1_mux_sel;
	wire input_addr_gen_1_restart;
	wire input_addr_gen_1_step;
	wire [7:0] output_addr_gen_0_addr_out;
	wire [2:0] output_addr_gen_0_mux_sel;
	wire output_addr_gen_0_restart;
	wire output_addr_gen_0_step;
	wire [7:0] output_addr_gen_1_addr_out;
	wire [2:0] output_addr_gen_1_mux_sel;
	wire output_addr_gen_1_restart;
	wire output_addr_gen_1_step;
	wire read;
	wire [31:0] s_read_addr;
	wire [31:0] s_write_addr;
	wire [31:0] sram_write_data;
	wire write;
	assign input_addr_gen_0_step = agg_read[0];
	assign input_addr_gen_0_restart = floop_restart[0];
	assign input_addr_gen_0_mux_sel = floop_mux_sel[0+:3];
	assign s_write_addr[7-:8] = input_addr_gen_0_addr_out;
	assign s_write_addr[15-:8] = 8'h00;
	assign input_addr_gen_1_step = agg_read[1];
	assign input_addr_gen_1_restart = floop_restart[1];
	assign input_addr_gen_1_mux_sel = floop_mux_sel[3+:3];
	assign s_write_addr[23-:8] = input_addr_gen_1_addr_out;
	assign s_write_addr[31-:8] = 8'h00;
	assign output_addr_gen_0_step = t_read[0];
	// assign output_addr_gen_0_restart = loops_sram2tb_restart[0];
	// assign output_addr_gen_0_mux_sel = loops_sram2tb_mux_sel[0+:3];
	assign s_read_addr[7-:8] = output_addr_gen_0_addr_out;
	assign s_read_addr[15-:8] = 8'h00;
	assign output_addr_gen_1_step = t_read[1];
	// assign output_addr_gen_1_restart = loops_sram2tb_restart[1];
	// assign output_addr_gen_1_mux_sel = loops_sram2tb_mux_sel[3+:3];

	// 给这些信号添加默认值
	assign output_addr_gen_0_mux_sel = 3'b0;
	assign output_addr_gen_0_restart = 1'b0;
	assign output_addr_gen_1_mux_sel = 3'b0;
	assign output_addr_gen_1_restart = 1'b0;

	assign s_read_addr[23-:8] = output_addr_gen_1_addr_out;
	assign s_read_addr[31-:8] = 8'h00;
	assign data_to_sram = sram_write_data;
	assign wen_to_sram = write;
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	always @(*) begin
		decode_sel_done_agg_read_s_write_addr = 1'h0;
		decode_ret_agg_read_s_write_addr = 16'h0000;
		begin : sv2v_autoblock_8
			reg [31:0] i;
			for (i = 0; i < 2; i = i + 1)
				if (~decode_sel_done_agg_read_s_write_addr & agg_read[sv2v_cast_1(i)]) begin
					decode_ret_agg_read_s_write_addr = s_write_addr[sv2v_cast_1(i) * 16+:16];
					decode_sel_done_agg_read_s_write_addr = 1'h1;
				end
		end
	end
	always @(*) begin
		decode_sel_done_t_read_s_read_addr = 1'h0;
		decode_ret_t_read_s_read_addr = 16'h0000;
		begin : sv2v_autoblock_9
			reg [31:0] i;
			for (i = 0; i < 2; i = i + 1)
				if (~decode_sel_done_t_read_s_read_addr & t_read[sv2v_cast_1(i)]) begin
					decode_ret_t_read_s_read_addr = s_read_addr[sv2v_cast_1(i) * 16+:16];
					decode_sel_done_t_read_s_read_addr = 1'h1;
				end
		end
	end
	assign ren_to_sram = read;
	assign wr_addr_to_sram = decode_ret_agg_read_s_write_addr[7:0];
	assign rd_addr_to_sram = decode_ret_t_read_s_read_addr[7:0];
	assign write = |agg_read;
	assign read = |t_read;
	always @(*) begin
		decode_sel_done_agg_read_agg_data_out = 1'h0;
		decode_ret_agg_read_agg_data_out = 32'h00000000;
		begin : sv2v_autoblock_10
			reg [31:0] i;
			for (i = 0; i < 2; i = i + 1)
				if (~decode_sel_done_agg_read_agg_data_out & agg_read[sv2v_cast_1(i)]) begin
					decode_ret_agg_read_agg_data_out = agg_data_out[16 * (sv2v_cast_1(i) * 2)+:32];
					decode_sel_done_agg_read_agg_data_out = 1'h1;
				end
		end
	end
	assign sram_write_data = decode_ret_agg_read_agg_data_out;
	addr_gen_6_8 input_addr_gen_0(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(input_addr_gen_0_mux_sel),
		.restart(input_addr_gen_0_restart),
		.rst_n(rst_n),
		.starting_addr(input_addr_gen_0_starting_addr),
		.step(input_addr_gen_0_step),
		.strides(input_addr_gen_0_strides),
		.addr_out(input_addr_gen_0_addr_out)
	);
	addr_gen_6_8 input_addr_gen_1(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(input_addr_gen_1_mux_sel),
		.restart(input_addr_gen_1_restart),
		.rst_n(rst_n),
		.starting_addr(input_addr_gen_1_starting_addr),
		.step(input_addr_gen_1_step),
		.strides(input_addr_gen_1_strides),
		.addr_out(input_addr_gen_1_addr_out)
	);
	addr_gen_6_8 output_addr_gen_0(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(output_addr_gen_0_mux_sel),
		.restart(output_addr_gen_0_restart),
		.rst_n(rst_n),
		.starting_addr(output_addr_gen_0_starting_addr),
		.step(output_addr_gen_0_step),
		.strides(output_addr_gen_0_strides),
		.addr_out(output_addr_gen_0_addr_out)
	);
	addr_gen_6_8 output_addr_gen_1(
		.clk(clk),
		.clk_en(clk_en),
		.flush(flush),
		.mux_sel(output_addr_gen_1_mux_sel),
		.restart(output_addr_gen_1_restart),
		.rst_n(rst_n),
		.starting_addr(output_addr_gen_1_starting_addr),
		.step(output_addr_gen_1_step),
		.strides(output_addr_gen_1_strides),
		.addr_out(output_addr_gen_1_addr_out)
	);
endmodule

// strg_ub_sram_tb_shared: 用于SRAM和测试模块之间的数据共享
// module strg_ub_sram_tb_shared (
// 	clk,
// 	clk_en,
// 	cycle_count,
// 	flush,
// 	loops_buf2out_autovec_read_0_dimensionality,
// 	loops_buf2out_autovec_read_0_ranges,
// 	loops_buf2out_autovec_read_1_dimensionality,
// 	loops_buf2out_autovec_read_1_ranges,
// 	output_sched_gen_0_enable,
// 	output_sched_gen_0_sched_addr_gen_starting_addr,
// 	output_sched_gen_0_sched_addr_gen_strides,
// 	output_sched_gen_1_enable,
// 	output_sched_gen_1_sched_addr_gen_starting_addr,
// 	output_sched_gen_1_sched_addr_gen_strides,
// 	rst_n,
// 	loops_sram2tb_mux_sel,
// 	loops_sram2tb_restart,
// 	t_read_out
// );
// 	input wire clk;
// 	input wire clk_en;
// 	input wire [15:0] cycle_count;
// 	input wire flush;
// 	input wire [3:0] loops_buf2out_autovec_read_0_dimensionality;
// 	input wire [95:0] loops_buf2out_autovec_read_0_ranges;
// 	input wire [3:0] loops_buf2out_autovec_read_1_dimensionality;
// 	input wire [95:0] loops_buf2out_autovec_read_1_ranges;
// 	input wire output_sched_gen_0_enable;
// 	input wire [15:0] output_sched_gen_0_sched_addr_gen_starting_addr;
// 	input wire [95:0] output_sched_gen_0_sched_addr_gen_strides;
// 	input wire output_sched_gen_1_enable;
// 	input wire [15:0] output_sched_gen_1_sched_addr_gen_starting_addr;
// 	input wire [95:0] output_sched_gen_1_sched_addr_gen_strides;
// 	input wire rst_n;
// 	output wire [5:0] loops_sram2tb_mux_sel;
// 	output wire [1:0] loops_sram2tb_restart;
// 	output wire [1:0] t_read_out;
// 	wire [2:0] loops_buf2out_autovec_read_0_mux_sel_out;
// 	wire loops_buf2out_autovec_read_0_restart;
// 	wire loops_buf2out_autovec_read_0_step;
// 	wire [2:0] loops_buf2out_autovec_read_1_mux_sel_out;
// 	wire loops_buf2out_autovec_read_1_restart;
// 	wire loops_buf2out_autovec_read_1_step;
// 	wire output_sched_gen_0_valid_output;
// 	wire output_sched_gen_1_valid_output;
// 	wire [1:0] t_read;
// 	assign t_read_out = t_read;
// 	assign loops_buf2out_autovec_read_0_step = t_read[0];
// 	assign loops_sram2tb_mux_sel[0+:3] = loops_buf2out_autovec_read_0_mux_sel_out;
// 	assign loops_sram2tb_restart[0] = loops_buf2out_autovec_read_0_restart;
// 	assign t_read[0] = output_sched_gen_0_valid_output;
// 	assign loops_buf2out_autovec_read_1_step = t_read[1];
// 	assign loops_sram2tb_mux_sel[3+:3] = loops_buf2out_autovec_read_1_mux_sel_out;
// 	assign loops_sram2tb_restart[1] = loops_buf2out_autovec_read_1_restart;
// 	assign t_read[1] = output_sched_gen_1_valid_output;
// 	for_loop_6_16 #(
// 		.CONFIG_WIDTH(5'h10),
// 		.ITERATOR_SUPPORT(4'h6)
// 	) loops_buf2out_autovec_read_0(
// 		.clk(clk),
// 		.clk_en(clk_en),
// 		.dimensionality(loops_buf2out_autovec_read_0_dimensionality),
// 		.flush(flush),
// 		.ranges(loops_buf2out_autovec_read_0_ranges),
// 		.rst_n(rst_n),
// 		.step(loops_buf2out_autovec_read_0_step),
// 		.mux_sel_out(loops_buf2out_autovec_read_0_mux_sel_out),
// 		.restart(loops_buf2out_autovec_read_0_restart)
// 	);
// 	sched_gen_6_16 output_sched_gen_0(
// 		.clk(clk),
// 		.clk_en(clk_en),
// 		.cycle_count(cycle_count),
// 		.enable(output_sched_gen_0_enable),
// 		.finished(loops_buf2out_autovec_read_0_restart),
// 		.flush(flush),
// 		.mux_sel(loops_buf2out_autovec_read_0_mux_sel_out),
// 		.rst_n(rst_n),
// 		.sched_addr_gen_starting_addr(output_sched_gen_0_sched_addr_gen_starting_addr),
// 		.sched_addr_gen_strides(output_sched_gen_0_sched_addr_gen_strides),
// 		.valid_output(output_sched_gen_0_valid_output)
// 	);
// 	for_loop_6_16 #(
// 		.CONFIG_WIDTH(5'h10),
// 		.ITERATOR_SUPPORT(4'h6)
// 	) loops_buf2out_autovec_read_1(
// 		.clk(clk),
// 		.clk_en(clk_en),
// 		.dimensionality(loops_buf2out_autovec_read_1_dimensionality),
// 		.flush(flush),
// 		.ranges(loops_buf2out_autovec_read_1_ranges),
// 		.rst_n(rst_n),
// 		.step(loops_buf2out_autovec_read_1_step),
// 		.mux_sel_out(loops_buf2out_autovec_read_1_mux_sel_out),
// 		.restart(loops_buf2out_autovec_read_1_restart)
// 	);
// 	sched_gen_6_16 output_sched_gen_1(
// 		.clk(clk),
// 		.clk_en(clk_en),
// 		.cycle_count(cycle_count),
// 		.enable(output_sched_gen_1_enable),
// 		.finished(loops_buf2out_autovec_read_1_restart),
// 		.flush(flush),
// 		.mux_sel(loops_buf2out_autovec_read_1_mux_sel_out),
// 		.rst_n(rst_n),
// 		.sched_addr_gen_starting_addr(output_sched_gen_1_sched_addr_gen_starting_addr),
// 		.sched_addr_gen_strides(output_sched_gen_1_sched_addr_gen_strides),
// 		.valid_output(output_sched_gen_1_valid_output)
// 	);
// endmodule

// strg_ub_tb_only: 模拟SRAM的读取行为，用于测试
// module strg_ub_tb_only (
// 	clk,
// 	clk_en,
// 	cycle_count,
// 	flush,
// 	loops_buf2out_read_0_dimensionality,
// 	loops_buf2out_read_0_ranges,
// 	loops_buf2out_read_1_dimensionality,
// 	loops_buf2out_read_1_ranges,
// 	loops_sram2tb_mux_sel,
// 	loops_sram2tb_restart,
// 	rst_n,
// 	sram_read_data,
// 	t_read,
// 	tb_read_addr_gen_0_starting_addr,
// 	tb_read_addr_gen_0_strides,
// 	tb_read_addr_gen_1_starting_addr,
// 	tb_read_addr_gen_1_strides,
// 	tb_read_sched_gen_0_enable,
// 	tb_read_sched_gen_0_sched_addr_gen_starting_addr,
// 	tb_read_sched_gen_0_sched_addr_gen_strides,
// 	tb_read_sched_gen_1_enable,
// 	tb_read_sched_gen_1_sched_addr_gen_starting_addr,
// 	tb_read_sched_gen_1_sched_addr_gen_strides,
// 	tb_write_addr_gen_0_starting_addr,
// 	tb_write_addr_gen_0_strides,
// 	tb_write_addr_gen_1_starting_addr,
// 	tb_write_addr_gen_1_strides,
// 	accessor_output,
// 	data_out
// );
// 	input wire clk;
// 	input wire clk_en;
// 	input wire [15:0] cycle_count;
// 	input wire flush;
// 	input wire [3:0] loops_buf2out_read_0_dimensionality;
// 	input wire [95:0] loops_buf2out_read_0_ranges;
// 	input wire [3:0] loops_buf2out_read_1_dimensionality;
// 	input wire [95:0] loops_buf2out_read_1_ranges;
// 	input wire [5:0] loops_sram2tb_mux_sel;
// 	input wire [1:0] loops_sram2tb_restart;
// 	input wire rst_n;
// 	input wire [31:0] sram_read_data;
// 	input wire [1:0] t_read;
// 	input wire [3:0] tb_read_addr_gen_0_starting_addr;
// 	input wire [23:0] tb_read_addr_gen_0_strides;
// 	input wire [3:0] tb_read_addr_gen_1_starting_addr;
// 	input wire [23:0] tb_read_addr_gen_1_strides;
// 	input wire tb_read_sched_gen_0_enable;
// 	input wire [15:0] tb_read_sched_gen_0_sched_addr_gen_starting_addr;
// 	input wire [95:0] tb_read_sched_gen_0_sched_addr_gen_strides;
// 	input wire tb_read_sched_gen_1_enable;
// 	input wire [15:0] tb_read_sched_gen_1_sched_addr_gen_starting_addr;
// 	input wire [95:0] tb_read_sched_gen_1_sched_addr_gen_strides;
// 	input wire [3:0] tb_write_addr_gen_0_starting_addr;
// 	input wire [23:0] tb_write_addr_gen_0_strides;
// 	input wire [3:0] tb_write_addr_gen_1_starting_addr;
// 	input wire [23:0] tb_write_addr_gen_1_strides;
// 	output wire [1:0] accessor_output;
// 	output reg [31:0] data_out;
// 	wire [2:0] loops_buf2out_read_0_mux_sel_out;
// 	wire loops_buf2out_read_0_restart;
// 	wire loops_buf2out_read_0_step;
// 	wire [2:0] loops_buf2out_read_1_mux_sel_out;
// 	wire loops_buf2out_read_1_restart;
// 	wire loops_buf2out_read_1_step;
// 	reg [5:0] mux_sel_d1;
// 	reg [1:0] restart_d1;
// 	reg [1:0] t_read_d1;
// 	reg [127:0] tb;
// 	wire [1:0] tb_read;
// 	wire [5:0] tb_read_addr;
// 	wire [3:0] tb_read_addr_gen_0_addr_out;
// 	wire tb_read_addr_gen_0_step;
// 	wire [3:0] tb_read_addr_gen_1_addr_out;
// 	wire tb_read_addr_gen_1_step;
// 	wire tb_read_sched_gen_0_valid_output;
// 	wire tb_read_sched_gen_1_valid_output;
// 	wire [5:0] tb_write_addr;
// 	wire [3:0] tb_write_addr_gen_0_addr_out;
// 	wire [2:0] tb_write_addr_gen_0_mux_sel;
// 	wire tb_write_addr_gen_0_restart;
// 	wire tb_write_addr_gen_0_step;
// 	wire [3:0] tb_write_addr_gen_1_addr_out;
// 	wire [2:0] tb_write_addr_gen_1_mux_sel;
// 	wire tb_write_addr_gen_1_restart;
// 	wire tb_write_addr_gen_1_step;
// 	assign accessor_output = tb_read;
// 	always @(posedge clk or negedge rst_n)
// 		if (~rst_n) begin
// 			t_read_d1[0] <= 1'h0;
// 			mux_sel_d1[0+:3] <= 3'h0;
// 			restart_d1[0] <= 1'h0;
// 		end
// 		else if (clk_en)
// 			if (flush) begin
// 				t_read_d1[0] <= 1'h0;
// 				mux_sel_d1[0+:3] <= 3'h0;
// 				restart_d1[0] <= 1'h0;
// 			end
// 			else begin
// 				t_read_d1[0] <= t_read[0];
// 				mux_sel_d1[0+:3] <= loops_sram2tb_mux_sel[0+:3];
// 				restart_d1[0] <= loops_sram2tb_restart[0];
// 			end
// 	always @(posedge clk or negedge rst_n)
// 		if (~rst_n) begin
// 			t_read_d1[1] <= 1'h0;
// 			mux_sel_d1[3+:3] <= 3'h0;
// 			restart_d1[1] <= 1'h0;
// 		end
// 		else if (clk_en)
// 			if (flush) begin
// 				t_read_d1[1] <= 1'h0;
// 				mux_sel_d1[3+:3] <= 3'h0;
// 				restart_d1[1] <= 1'h0;
// 			end
// 			else begin
// 				t_read_d1[1] <= t_read[1];
// 				mux_sel_d1[3+:3] <= loops_sram2tb_mux_sel[3+:3];
// 				restart_d1[1] <= loops_sram2tb_restart[1];
// 			end
// 	assign tb_write_addr_gen_0_step = t_read_d1[0];
// 	assign tb_write_addr_gen_0_mux_sel = mux_sel_d1[0+:3];
// 	assign tb_write_addr_gen_0_restart = restart_d1[0];
// 	assign tb_write_addr[0+:3] = tb_write_addr_gen_0_addr_out[2:0];
// 	always @(posedge clk)
// 		if (clk_en)
// 			if (t_read_d1[0])
// 				tb[16 * (tb_write_addr[0] * 2)+:32] <= sram_read_data;
// 	assign loops_buf2out_read_0_step = tb_read[0];
// 	assign tb_read_addr_gen_0_step = tb_read[0];
// 	assign tb_read_addr[0+:3] = tb_read_addr_gen_0_addr_out[2:0];
// 	assign tb_read[0] = tb_read_sched_gen_0_valid_output;
// 	always @(*) data_out[0+:16] = tb[((tb_read_addr[1] * 2) + tb_read_addr[0]) * 16+:16];
// 	assign tb_write_addr_gen_1_step = t_read_d1[1];
// 	assign tb_write_addr_gen_1_mux_sel = mux_sel_d1[3+:3];
// 	assign tb_write_addr_gen_1_restart = restart_d1[1];
// 	assign tb_write_addr[3+:3] = tb_write_addr_gen_1_addr_out[2:0];
// 	always @(posedge clk)
// 		if (clk_en)
// 			if (t_read_d1[1])
// 				tb[16 * ((2 + tb_write_addr[3]) * 2)+:32] <= sram_read_data;
// 	assign loops_buf2out_read_1_step = tb_read[1];
// 	assign tb_read_addr_gen_1_step = tb_read[1];
// 	assign tb_read_addr[3+:3] = tb_read_addr_gen_1_addr_out[2:0];
// 	assign tb_read[1] = tb_read_sched_gen_1_valid_output;
// 	always @(*) data_out[16+:16] = tb[(((2 + tb_read_addr[4]) * 2) + tb_read_addr[3]) * 16+:16];
// 	addr_gen_6_4 tb_write_addr_gen_0(
// 		.clk(clk),
// 		.clk_en(clk_en),
// 		.flush(flush),
// 		.mux_sel(tb_write_addr_gen_0_mux_sel),
// 		.restart(tb_write_addr_gen_0_restart),
// 		.rst_n(rst_n),
// 		.starting_addr(tb_write_addr_gen_0_starting_addr),
// 		.step(tb_write_addr_gen_0_step),
// 		.strides(tb_write_addr_gen_0_strides),
// 		.addr_out(tb_write_addr_gen_0_addr_out)
// 	);
// 	for_loop_6_16 #(
// 		.CONFIG_WIDTH(5'h10),
// 		.ITERATOR_SUPPORT(4'h6)
// 	) loops_buf2out_read_0(
// 		.clk(clk),
// 		.clk_en(clk_en),
// 		.dimensionality(loops_buf2out_read_0_dimensionality),
// 		.flush(flush),
// 		.ranges(loops_buf2out_read_0_ranges),
// 		.rst_n(rst_n),
// 		.step(loops_buf2out_read_0_step),
// 		.mux_sel_out(loops_buf2out_read_0_mux_sel_out),
// 		.restart(loops_buf2out_read_0_restart)
// 	);
// 	addr_gen_6_4 tb_read_addr_gen_0(
// 		.clk(clk),
// 		.clk_en(clk_en),
// 		.flush(flush),
// 		.mux_sel(loops_buf2out_read_0_mux_sel_out),
// 		.restart(loops_buf2out_read_0_restart),
// 		.rst_n(rst_n),
// 		.starting_addr(tb_read_addr_gen_0_starting_addr),
// 		.step(tb_read_addr_gen_0_step),
// 		.strides(tb_read_addr_gen_0_strides),
// 		.addr_out(tb_read_addr_gen_0_addr_out)
// 	);
// 	sched_gen_6_16 tb_read_sched_gen_0(
// 		.clk(clk),
// 		.clk_en(clk_en),
// 		.cycle_count(cycle_count),
// 		.enable(tb_read_sched_gen_0_enable),
// 		.finished(loops_buf2out_read_0_restart),
// 		.flush(flush),
// 		.mux_sel(loops_buf2out_read_0_mux_sel_out),
// 		.rst_n(rst_n),
// 		.sched_addr_gen_starting_addr(tb_read_sched_gen_0_sched_addr_gen_starting_addr),
// 		.sched_addr_gen_strides(tb_read_sched_gen_0_sched_addr_gen_strides),
// 		.valid_output(tb_read_sched_gen_0_valid_output)
// 	);
// 	addr_gen_6_4 tb_write_addr_gen_1(
// 		.clk(clk),
// 		.clk_en(clk_en),
// 		.flush(flush),
// 		.mux_sel(tb_write_addr_gen_1_mux_sel),
// 		.restart(tb_write_addr_gen_1_restart),
// 		.rst_n(rst_n),
// 		.starting_addr(tb_write_addr_gen_1_starting_addr),
// 		.step(tb_write_addr_gen_1_step),
// 		.strides(tb_write_addr_gen_1_strides),
// 		.addr_out(tb_write_addr_gen_1_addr_out)
// 	);
// 	for_loop_6_16 #(
// 		.CONFIG_WIDTH(5'h10),
// 		.ITERATOR_SUPPORT(4'h6)
// 	) loops_buf2out_read_1(
// 		.clk(clk),
// 		.clk_en(clk_en),
// 		.dimensionality(loops_buf2out_read_1_dimensionality),
// 		.flush(flush),
// 		.ranges(loops_buf2out_read_1_ranges),
// 		.rst_n(rst_n),
// 		.step(loops_buf2out_read_1_step),
// 		.mux_sel_out(loops_buf2out_read_1_mux_sel_out),
// 		.restart(loops_buf2out_read_1_restart)
// 	);
// 	addr_gen_6_4 tb_read_addr_gen_1(
// 		.clk(clk),
// 		.clk_en(clk_en),
// 		.flush(flush),
// 		.mux_sel(loops_buf2out_read_1_mux_sel_out),
// 		.restart(loops_buf2out_read_1_restart),
// 		.rst_n(rst_n),
// 		.starting_addr(tb_read_addr_gen_1_starting_addr),
// 		.step(tb_read_addr_gen_1_step),
// 		.strides(tb_read_addr_gen_1_strides),
// 		.addr_out(tb_read_addr_gen_1_addr_out)
// 	);
// 	sched_gen_6_16 tb_read_sched_gen_1(
// 		.clk(clk),
// 		.clk_en(clk_en),
// 		.cycle_count(cycle_count),
// 		.enable(tb_read_sched_gen_1_enable),
// 		.finished(loops_buf2out_read_1_restart),
// 		.flush(flush),
// 		.mux_sel(loops_buf2out_read_1_mux_sel_out),
// 		.rst_n(rst_n),
// 		.sched_addr_gen_starting_addr(tb_read_sched_gen_1_sched_addr_gen_starting_addr),
// 		.sched_addr_gen_strides(tb_read_sched_gen_1_sched_addr_gen_strides),
// 		.valid_output(tb_read_sched_gen_1_valid_output)
// 	);
// endmodule
module strg_ub_vec (
	agg_only_agg_read_addr_gen_0_starting_addr,
	agg_only_agg_read_addr_gen_0_strides,
	agg_only_agg_read_addr_gen_1_starting_addr,
	agg_only_agg_read_addr_gen_1_strides,
	agg_only_agg_write_addr_gen_0_starting_addr,
	agg_only_agg_write_addr_gen_0_strides,
	agg_only_agg_write_addr_gen_1_starting_addr,
	agg_only_agg_write_addr_gen_1_strides,
	agg_only_agg_write_sched_gen_0_enable,
	agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr,
	agg_only_agg_write_sched_gen_0_sched_addr_gen_strides,
	agg_only_agg_write_sched_gen_1_enable,
	agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr,
	agg_only_agg_write_sched_gen_1_sched_addr_gen_strides,
	agg_only_loops_in2buf_0_dimensionality,
	agg_only_loops_in2buf_0_ranges,
	agg_only_loops_in2buf_1_dimensionality,
	agg_only_loops_in2buf_1_ranges,
	agg_sram_shared_agg_read_sched_gen_0_enable,
	agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr,
	agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides,
	agg_sram_shared_agg_read_sched_gen_1_enable,
	agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr,
	agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides,
	agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality,
	agg_sram_shared_loops_in2buf_autovec_write_0_ranges,
	agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality,
	agg_sram_shared_loops_in2buf_autovec_write_1_ranges,
	chain_chain_en,
	chain_data_in,
	clk,
	clk_en,
	data_from_strg,
	data_in,
	flush,
	rst_n,
	sram_only_input_addr_gen_0_starting_addr,
	sram_only_input_addr_gen_0_strides,
	sram_only_input_addr_gen_1_starting_addr,
	sram_only_input_addr_gen_1_strides,
	sram_only_output_addr_gen_0_starting_addr,
	sram_only_output_addr_gen_0_strides,
	sram_only_output_addr_gen_1_starting_addr,
	sram_only_output_addr_gen_1_strides,
	// sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality,
	// sram_tb_shared_loops_buf2out_autovec_read_0_ranges,
	// sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality,
	// sram_tb_shared_loops_buf2out_autovec_read_1_ranges,
	// sram_tb_shared_output_sched_gen_0_enable,
	// sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr,
	// sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides,
	// sram_tb_shared_output_sched_gen_1_enable,
	// sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr,
	// sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides,
	// tb_only_loops_buf2out_read_0_dimensionality,
	// tb_only_loops_buf2out_read_0_ranges,
	// tb_only_loops_buf2out_read_1_dimensionality,
	// tb_only_loops_buf2out_read_1_ranges,
	// tb_only_tb_read_addr_gen_0_starting_addr,
	// tb_only_tb_read_addr_gen_0_strides,
	// tb_only_tb_read_addr_gen_1_starting_addr,
	// tb_only_tb_read_addr_gen_1_strides,
	// tb_only_tb_read_sched_gen_0_enable,
	// tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr,
	// tb_only_tb_read_sched_gen_0_sched_addr_gen_strides,
	// tb_only_tb_read_sched_gen_1_enable,
	// tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr,
	// tb_only_tb_read_sched_gen_1_sched_addr_gen_strides,
	// tb_only_tb_write_addr_gen_0_starting_addr,
	// tb_only_tb_write_addr_gen_0_strides,
	// tb_only_tb_write_addr_gen_1_starting_addr,
	// tb_only_tb_write_addr_gen_1_strides,
	accessor_output,
	data_out,
	data_to_strg,
	rd_addr_out,
	ren_to_strg,
	tmp0_rdaddr,
	tmp0_rden,
	wen_to_strg,
	wr_addr_out
);
	input wire [3:0] agg_only_agg_read_addr_gen_0_starting_addr;
	input wire [23:0] agg_only_agg_read_addr_gen_0_strides;
	input wire [3:0] agg_only_agg_read_addr_gen_1_starting_addr;
	input wire [23:0] agg_only_agg_read_addr_gen_1_strides;
	input wire [3:0] agg_only_agg_write_addr_gen_0_starting_addr;
	input wire [23:0] agg_only_agg_write_addr_gen_0_strides;
	input wire [3:0] agg_only_agg_write_addr_gen_1_starting_addr;
	input wire [23:0] agg_only_agg_write_addr_gen_1_strides;
	input wire agg_only_agg_write_sched_gen_0_enable;
	input wire [15:0] agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr;
	input wire [95:0] agg_only_agg_write_sched_gen_0_sched_addr_gen_strides;
	input wire agg_only_agg_write_sched_gen_1_enable;
	input wire [15:0] agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr;
	input wire [95:0] agg_only_agg_write_sched_gen_1_sched_addr_gen_strides;
	input wire [3:0] agg_only_loops_in2buf_0_dimensionality;
	input wire [95:0] agg_only_loops_in2buf_0_ranges;
	input wire [3:0] agg_only_loops_in2buf_1_dimensionality;
	input wire [95:0] agg_only_loops_in2buf_1_ranges;
	input wire agg_sram_shared_agg_read_sched_gen_0_enable;
	input wire [15:0] agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr;
	input wire [95:0] agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides;
	input wire agg_sram_shared_agg_read_sched_gen_1_enable;
	input wire [15:0] agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr;
	input wire [95:0] agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides;
	input wire [3:0] agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality;
	input wire [95:0] agg_sram_shared_loops_in2buf_autovec_write_0_ranges;
	input wire [3:0] agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality;
	input wire [95:0] agg_sram_shared_loops_in2buf_autovec_write_1_ranges;
	input wire chain_chain_en;
	input wire [31:0] chain_data_in;
	input wire clk;
	input wire clk_en;
	input wire [31:0] data_from_strg; // 来自 SRAM 的数据
	input wire [31:0] data_in;
	input wire flush;
	input wire rst_n;
	input wire [7:0] sram_only_input_addr_gen_0_starting_addr;
	input wire [47:0] sram_only_input_addr_gen_0_strides;
	input wire [7:0] sram_only_input_addr_gen_1_starting_addr;
	input wire [47:0] sram_only_input_addr_gen_1_strides;
	input wire [7:0] sram_only_output_addr_gen_0_starting_addr;
	input wire [47:0] sram_only_output_addr_gen_0_strides;
	input wire [7:0] sram_only_output_addr_gen_1_starting_addr;
	input wire [47:0] sram_only_output_addr_gen_1_strides;
	// input wire [3:0] sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality;
	// input wire [95:0] sram_tb_shared_loops_buf2out_autovec_read_0_ranges;
	// input wire [3:0] sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality;
	// input wire [95:0] sram_tb_shared_loops_buf2out_autovec_read_1_ranges;
	// input wire sram_tb_shared_output_sched_gen_0_enable;
	// input wire [15:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr;
	// input wire [95:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides;
	// input wire sram_tb_shared_output_sched_gen_1_enable;
	// input wire [15:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr;
	// input wire [95:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides;
	// input wire [3:0] tb_only_loops_buf2out_read_0_dimensionality;
	// input wire [95:0] tb_only_loops_buf2out_read_0_ranges;
	// input wire [3:0] tb_only_loops_buf2out_read_1_dimensionality;
	// input wire [95:0] tb_only_loops_buf2out_read_1_ranges;
	// input wire [3:0] tb_only_tb_read_addr_gen_0_starting_addr;
	// input wire [23:0] tb_only_tb_read_addr_gen_0_strides;
	// input wire [3:0] tb_only_tb_read_addr_gen_1_starting_addr;
	// input wire [23:0] tb_only_tb_read_addr_gen_1_strides;
	// input wire tb_only_tb_read_sched_gen_0_enable;
	// input wire [15:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr;
	// input wire [95:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_strides;
	// input wire tb_only_tb_read_sched_gen_1_enable;
	// input wire [15:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr;
	// input wire [95:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_strides;
	// input wire [3:0] tb_only_tb_write_addr_gen_0_starting_addr;
	// input wire [23:0] tb_only_tb_write_addr_gen_0_strides;
	// input wire [3:0] tb_only_tb_write_addr_gen_1_starting_addr;
	// input wire [23:0] tb_only_tb_write_addr_gen_1_strides;
	output wire [1:0] accessor_output;
	output wire [31:0] data_out; // 输出到 Tile 的数据
	output wire [31:0] data_to_strg; // 给 SRAM 的数据
	output wire [7:0] rd_addr_out;
	output wire ren_to_strg;
	output wire [7:0] tmp0_rdaddr;
	output wire tmp0_rden;
	output wire wen_to_strg;
	output wire [7:0] wr_addr_out;
	wire [1:0] accessor_output_int; // 只连接到了strg_ub_tb_only 模块, 没有实际的驱动源
	wire [63:0] agg_only_agg_data_out;
	wire [1:0] agg_only_agg_read;
	wire [5:0] agg_only_floop_mux_sel;
	wire [1:0] agg_only_floop_restart;
	wire [1:0] agg_sram_shared_agg_read_out;
	wire [5:0] agg_sram_shared_floop_mux_sel;
	wire [1:0] agg_sram_shared_floop_restart;
	reg [15:0] cycle_count;
	wire [31:0] data_out_int; // 这个信号是 strg_ub_tb_only 模块的输入，在 RTL 代码中没有驱动源
	// wire [5:0] sram_only_loops_sram2tb_mux_sel;
	// wire [1:0] sram_only_loops_sram2tb_restart;
	// wire [1:0] sram_only_t_read; // 这个信号只连接到了 strg_ub_tb_only 模块
	// wire [5:0] sram_tb_shared_loops_sram2tb_mux_sel;
	// wire [1:0] sram_tb_shared_loops_sram2tb_restart;
	// wire [1:0] sram_tb_shared_t_read_out;
	always @(posedge clk or negedge rst_n)
		if (~rst_n)
			cycle_count <= 16'h0000;
		else if (clk_en)
			if (flush)
				cycle_count <= 16'h0000;
			else
				cycle_count <= cycle_count + 16'h0001;
	assign agg_only_agg_read = agg_sram_shared_agg_read_out;
	assign agg_only_floop_mux_sel = agg_sram_shared_floop_mux_sel;
	assign agg_only_floop_restart = agg_sram_shared_floop_restart;
	// assign sram_only_loops_sram2tb_mux_sel = sram_tb_shared_loops_sram2tb_mux_sel;
	// assign sram_only_loops_sram2tb_restart = sram_tb_shared_loops_sram2tb_restart;
	// assign sram_only_t_read = sram_tb_shared_t_read_out;
	assign tmp0_rdaddr = 8'h00;
	assign tmp0_rden = 1'h0;
	assign accessor_output = accessor_output_int;
	strg_ub_agg_only agg_only(
		.agg_read(agg_only_agg_read),
		.agg_read_addr_gen_0_starting_addr(agg_only_agg_read_addr_gen_0_starting_addr),
		.agg_read_addr_gen_0_strides(agg_only_agg_read_addr_gen_0_strides),
		.agg_read_addr_gen_1_starting_addr(agg_only_agg_read_addr_gen_1_starting_addr),
		.agg_read_addr_gen_1_strides(agg_only_agg_read_addr_gen_1_strides),
		.agg_write_addr_gen_0_starting_addr(agg_only_agg_write_addr_gen_0_starting_addr),
		.agg_write_addr_gen_0_strides(agg_only_agg_write_addr_gen_0_strides),
		.agg_write_addr_gen_1_starting_addr(agg_only_agg_write_addr_gen_1_starting_addr),
		.agg_write_addr_gen_1_strides(agg_only_agg_write_addr_gen_1_strides),
		.agg_write_sched_gen_0_enable(agg_only_agg_write_sched_gen_0_enable),
		.agg_write_sched_gen_0_sched_addr_gen_starting_addr(agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr),
		.agg_write_sched_gen_0_sched_addr_gen_strides(agg_only_agg_write_sched_gen_0_sched_addr_gen_strides),
		.agg_write_sched_gen_1_enable(agg_only_agg_write_sched_gen_1_enable),
		.agg_write_sched_gen_1_sched_addr_gen_starting_addr(agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr),
		.agg_write_sched_gen_1_sched_addr_gen_strides(agg_only_agg_write_sched_gen_1_sched_addr_gen_strides),
		.clk(clk),
		.clk_en(clk_en),
		.cycle_count(cycle_count),
		.data_in(data_in),
		.floop_mux_sel(agg_only_floop_mux_sel),
		.floop_restart(agg_only_floop_restart),
		.flush(flush),
		.loops_in2buf_0_dimensionality(agg_only_loops_in2buf_0_dimensionality),
		.loops_in2buf_0_ranges(agg_only_loops_in2buf_0_ranges),
		.loops_in2buf_1_dimensionality(agg_only_loops_in2buf_1_dimensionality),
		.loops_in2buf_1_ranges(agg_only_loops_in2buf_1_ranges),
		.rst_n(rst_n),
		.agg_data_out(agg_only_agg_data_out)
	);
	strg_ub_agg_sram_shared agg_sram_shared(
		.agg_read_sched_gen_0_enable(agg_sram_shared_agg_read_sched_gen_0_enable),
		.agg_read_sched_gen_0_sched_addr_gen_starting_addr(agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr),
		.agg_read_sched_gen_0_sched_addr_gen_strides(agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides),
		.agg_read_sched_gen_1_enable(agg_sram_shared_agg_read_sched_gen_1_enable),
		.agg_read_sched_gen_1_sched_addr_gen_starting_addr(agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr),
		.agg_read_sched_gen_1_sched_addr_gen_strides(agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides),
		.clk(clk),
		.clk_en(clk_en),
		.cycle_count(cycle_count),
		.flush(flush),
		.loops_in2buf_autovec_write_0_dimensionality(agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality),
		.loops_in2buf_autovec_write_0_ranges(agg_sram_shared_loops_in2buf_autovec_write_0_ranges),
		.loops_in2buf_autovec_write_1_dimensionality(agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality),
		.loops_in2buf_autovec_write_1_ranges(agg_sram_shared_loops_in2buf_autovec_write_1_ranges),
		.rst_n(rst_n),
		.agg_read_out(agg_sram_shared_agg_read_out),
		.floop_mux_sel(agg_sram_shared_floop_mux_sel),
		.floop_restart(agg_sram_shared_floop_restart)
	);
	strg_ub_sram_only sram_only(
		.agg_data_out(agg_only_agg_data_out),
		.agg_read(agg_sram_shared_agg_read_out),
		.clk(clk),
		.clk_en(clk_en),
		.cycle_count(cycle_count),
		.floop_mux_sel(agg_sram_shared_floop_mux_sel),
		.floop_restart(agg_sram_shared_floop_restart),
		.flush(flush),
		.input_addr_gen_0_starting_addr(sram_only_input_addr_gen_0_starting_addr),
		.input_addr_gen_0_strides(sram_only_input_addr_gen_0_strides),
		.input_addr_gen_1_starting_addr(sram_only_input_addr_gen_1_starting_addr),
		.input_addr_gen_1_strides(sram_only_input_addr_gen_1_strides),
		// .loops_sram2tb_mux_sel(sram_only_loops_sram2tb_mux_sel),
		// .loops_sram2tb_restart(sram_only_loops_sram2tb_restart),
		.output_addr_gen_0_starting_addr(sram_only_output_addr_gen_0_starting_addr),
		.output_addr_gen_0_strides(sram_only_output_addr_gen_0_strides),
		.output_addr_gen_1_starting_addr(sram_only_output_addr_gen_1_starting_addr),
		.output_addr_gen_1_strides(sram_only_output_addr_gen_1_strides),
		.rst_n(rst_n),
		// .t_read(sram_only_t_read),
		.data_to_sram(data_to_strg),
		.rd_addr_to_sram(rd_addr_out),
		.ren_to_sram(ren_to_strg),
		.wen_to_sram(wen_to_strg),
		.wr_addr_to_sram(wr_addr_out)
	);

	// strg_ub_sram_tb_shared: 用于SRAM和测试模块之间的数据共享
	// strg_ub_sram_tb_shared sram_tb_shared(
	// 	.clk(clk),
	// 	.clk_en(clk_en),
	// 	.cycle_count(cycle_count),
	// 	.flush(flush),
	// 	.loops_buf2out_autovec_read_0_dimensionality(sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality),
	// 	.loops_buf2out_autovec_read_0_ranges(sram_tb_shared_loops_buf2out_autovec_read_0_ranges),
	// 	.loops_buf2out_autovec_read_1_dimensionality(sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality),
	// 	.loops_buf2out_autovec_read_1_ranges(sram_tb_shared_loops_buf2out_autovec_read_1_ranges),
	// 	.output_sched_gen_0_enable(sram_tb_shared_output_sched_gen_0_enable),
	// 	.output_sched_gen_0_sched_addr_gen_starting_addr(sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr),
	// 	.output_sched_gen_0_sched_addr_gen_strides(sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides),
	// 	.output_sched_gen_1_enable(sram_tb_shared_output_sched_gen_1_enable),
	// 	.output_sched_gen_1_sched_addr_gen_starting_addr(sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr),
	// 	.output_sched_gen_1_sched_addr_gen_strides(sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides),
	// 	.rst_n(rst_n),
	// 	.loops_sram2tb_mux_sel(sram_tb_shared_loops_sram2tb_mux_sel),
	// 	.loops_sram2tb_restart(sram_tb_shared_loops_sram2tb_restart),
	// 	.t_read_out(sram_tb_shared_t_read_out)
	// );

	// strg_ub_tb_only: 模拟SRAM的读取行为，用于测试
	// strg_ub_tb_only tb_only(
	// 	.clk(clk),
	// 	.clk_en(clk_en),
	// 	.cycle_count(cycle_count),
	// 	.flush(flush),
	// 	.loops_buf2out_read_0_dimensionality(tb_only_loops_buf2out_read_0_dimensionality),
	// 	.loops_buf2out_read_0_ranges(tb_only_loops_buf2out_read_0_ranges),
	// 	.loops_buf2out_read_1_dimensionality(tb_only_loops_buf2out_read_1_dimensionality),
	// 	.loops_buf2out_read_1_ranges(tb_only_loops_buf2out_read_1_ranges),
	// 	.loops_sram2tb_mux_sel(sram_tb_shared_loops_sram2tb_mux_sel),
	// 	.loops_sram2tb_restart(sram_tb_shared_loops_sram2tb_restart),
	// 	.rst_n(rst_n),
	// 	.sram_read_data(data_from_strg),
	// 	.t_read(sram_tb_shared_t_read_out),
	// 	.tb_read_addr_gen_0_starting_addr(tb_only_tb_read_addr_gen_0_starting_addr),
	// 	.tb_read_addr_gen_0_strides(tb_only_tb_read_addr_gen_0_strides),
	// 	.tb_read_addr_gen_1_starting_addr(tb_only_tb_read_addr_gen_1_starting_addr),
	// 	.tb_read_addr_gen_1_strides(tb_only_tb_read_addr_gen_1_strides),
	// 	.tb_read_sched_gen_0_enable(tb_only_tb_read_sched_gen_0_enable),
	// 	.tb_read_sched_gen_0_sched_addr_gen_starting_addr(tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr),
	// 	.tb_read_sched_gen_0_sched_addr_gen_strides(tb_only_tb_read_sched_gen_0_sched_addr_gen_strides),
	// 	.tb_read_sched_gen_1_enable(tb_only_tb_read_sched_gen_1_enable),
	// 	.tb_read_sched_gen_1_sched_addr_gen_starting_addr(tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr),
	// 	.tb_read_sched_gen_1_sched_addr_gen_strides(tb_only_tb_read_sched_gen_1_sched_addr_gen_strides),
	// 	.tb_write_addr_gen_0_starting_addr(tb_only_tb_write_addr_gen_0_starting_addr),
	// 	.tb_write_addr_gen_0_strides(tb_only_tb_write_addr_gen_0_strides),
	// 	.tb_write_addr_gen_1_starting_addr(tb_only_tb_write_addr_gen_1_starting_addr),
	// 	.tb_write_addr_gen_1_strides(tb_only_tb_write_addr_gen_1_strides),
	// 	.accessor_output(accessor_output_int),
	// 	.data_out(data_out_int)
	// );

	// 屏蔽TestBench后，从SRAM部分获取数据
	assign data_out_int = data_from_strg;  // 假设data_from_strg是从SRAM读出的数据
	assign accessor_output_int = 2'b0;     // 需要根据实际需求设置适当的值

	Chain chain(
		.accessor_output(accessor_output_int),
		.chain_data_in(chain_data_in),
		.chain_en(chain_chain_en),
		.clk_en(clk_en),
		.curr_tile_data_out(data_out_int),
		.flush(flush),
		.data_out_tile(data_out)
	);
endmodule
module strg_ub_vec_flat (
	chain_data_in_f_0,
	chain_data_in_f_1,
	clk,
	clk_en,
	data_from_strg_lifted,
	data_in_f_0,
	data_in_f_1,
	flush,
	rst_n,
	strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr,
	strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides,
	strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr,
	strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides,
	strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr,
	strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides,
	strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr,
	strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides,
	strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable,
	strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr,
	strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides,
	strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable,
	strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr,
	strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides,
	strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality,
	strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges,
	strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality,
	strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges,
	strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable,
	strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr,
	strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides,
	strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable,
	strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr,
	strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides,
	strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality,
	strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges,
	strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality,
	strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges,
	strg_ub_vec_inst_chain_chain_en,
	strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr,
	strg_ub_vec_inst_sram_only_input_addr_gen_0_strides,
	strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr,
	strg_ub_vec_inst_sram_only_input_addr_gen_1_strides,
	strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr,
	strg_ub_vec_inst_sram_only_output_addr_gen_0_strides,
	strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr,
	strg_ub_vec_inst_sram_only_output_addr_gen_1_strides,
	// strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality,
	// strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges,
	// strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality,
	// strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges,
	// strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable,
	// strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr,
	// strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides,
	// strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable,
	// strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr,
	// strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides,
	// strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality,
	// strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges,
	// strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality,
	// strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges,
	// strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr,
	// strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides,
	// strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr,
	// strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides,
	// strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable,
	// strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr,
	// strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides,
	// strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable,
	// strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr,
	// strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides,
	// strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr,
	// strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides,
	// strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr,
	// strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides,
	accessor_output_f_b_0,
	accessor_output_f_b_1,
	data_out_f_0,
	data_out_f_1,
	data_to_strg_lifted,
	rd_addr_out_lifted,
	ren_to_strg_lifted,
	tmp0_rdaddr_lifted,
	tmp0_rden_lifted,
	wen_to_strg_lifted,
	wr_addr_out_lifted
);
	input wire [15:0] chain_data_in_f_0;
	input wire [15:0] chain_data_in_f_1;
	input wire clk;
	input wire clk_en;
	input wire [31:0] data_from_strg_lifted;
	input wire [15:0] data_in_f_0;
	input wire [15:0] data_in_f_1;
	input wire flush;
	input wire rst_n;
	input wire [3:0] strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr;
	input wire [23:0] strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides;
	input wire [3:0] strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr;
	input wire [23:0] strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides;
	input wire [3:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr;
	input wire [23:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides;
	input wire [3:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr;
	input wire [23:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides;
	input wire strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable;
	input wire [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr;
	input wire [95:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides;
	input wire strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable;
	input wire [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr;
	input wire [95:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides;
	input wire [3:0] strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality;
	input wire [95:0] strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges;
	input wire [3:0] strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality;
	input wire [95:0] strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges;
	input wire strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable;
	input wire [15:0] strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr;
	input wire [95:0] strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides;
	input wire strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable;
	input wire [15:0] strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr;
	input wire [95:0] strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides;
	input wire [3:0] strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality;
	input wire [95:0] strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges;
	input wire [3:0] strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality;
	input wire [95:0] strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges;
	input wire strg_ub_vec_inst_chain_chain_en;
	input wire [7:0] strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr;
	input wire [47:0] strg_ub_vec_inst_sram_only_input_addr_gen_0_strides;
	input wire [7:0] strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr;
	input wire [47:0] strg_ub_vec_inst_sram_only_input_addr_gen_1_strides;
	input wire [7:0] strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr;
	input wire [47:0] strg_ub_vec_inst_sram_only_output_addr_gen_0_strides;
	input wire [7:0] strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr;
	input wire [47:0] strg_ub_vec_inst_sram_only_output_addr_gen_1_strides;
	// input wire [3:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality;
	// input wire [95:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges;
	// input wire [3:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality;
	// input wire [95:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges;
	// input wire strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable;
	// input wire [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr;
	// input wire [95:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides;
	// input wire strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable;
	// input wire [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr;
	// input wire [95:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides;
	// input wire [3:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality;
	// input wire [95:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges;
	// input wire [3:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality;
	// input wire [95:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges;
	// input wire [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr;
	// input wire [23:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides;
	// input wire [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr;
	// input wire [23:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides;
	// input wire strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable;
	// input wire [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr;
	// input wire [95:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides;
	// input wire strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable;
	// input wire [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr;
	// input wire [95:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides;
	// input wire [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr;
	// input wire [23:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides;
	// input wire [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr;
	// input wire [23:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides;
	output wire accessor_output_f_b_0;
	output wire accessor_output_f_b_1;
	output wire [15:0] data_out_f_0;
	output wire [15:0] data_out_f_1;
	output wire [31:0] data_to_strg_lifted;
	output wire [7:0] rd_addr_out_lifted;
	output wire ren_to_strg_lifted;
	output wire [7:0] tmp0_rdaddr_lifted;
	output wire tmp0_rden_lifted;
	output wire wen_to_strg_lifted;
	output wire [7:0] wr_addr_out_lifted;
	wire [1:0] strg_ub_vec_inst_accessor_output;
	wire [31:0] strg_ub_vec_inst_chain_data_in;
	wire [31:0] strg_ub_vec_inst_data_in;
	wire [31:0] strg_ub_vec_inst_data_out;
	assign strg_ub_vec_inst_chain_data_in[0+:16] = chain_data_in_f_0;
	assign strg_ub_vec_inst_chain_data_in[16+:16] = chain_data_in_f_1;
	assign strg_ub_vec_inst_data_in[0+:16] = data_in_f_0;
	assign strg_ub_vec_inst_data_in[16+:16] = data_in_f_1;
	assign accessor_output_f_b_0 = strg_ub_vec_inst_accessor_output[0];
	assign accessor_output_f_b_1 = strg_ub_vec_inst_accessor_output[1];
	assign data_out_f_0 = strg_ub_vec_inst_data_out[0+:16];
	assign data_out_f_1 = strg_ub_vec_inst_data_out[16+:16];
	strg_ub_vec strg_ub_vec_inst(
		.agg_only_agg_read_addr_gen_0_starting_addr(strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr),
		.agg_only_agg_read_addr_gen_0_strides(strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides),
		.agg_only_agg_read_addr_gen_1_starting_addr(strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr),
		.agg_only_agg_read_addr_gen_1_strides(strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides),
		.agg_only_agg_write_addr_gen_0_starting_addr(strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr),
		.agg_only_agg_write_addr_gen_0_strides(strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides),
		.agg_only_agg_write_addr_gen_1_starting_addr(strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr),
		.agg_only_agg_write_addr_gen_1_strides(strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides),
		.agg_only_agg_write_sched_gen_0_enable(strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable),
		.agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr),
		.agg_only_agg_write_sched_gen_0_sched_addr_gen_strides(strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides),
		.agg_only_agg_write_sched_gen_1_enable(strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable),
		.agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr),
		.agg_only_agg_write_sched_gen_1_sched_addr_gen_strides(strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides),
		.agg_only_loops_in2buf_0_dimensionality(strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality),
		.agg_only_loops_in2buf_0_ranges(strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges),
		.agg_only_loops_in2buf_1_dimensionality(strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality),
		.agg_only_loops_in2buf_1_ranges(strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges),
		.agg_sram_shared_agg_read_sched_gen_0_enable(strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable),
		.agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr),
		.agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides(strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides),
		.agg_sram_shared_agg_read_sched_gen_1_enable(strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable),
		.agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr),
		.agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides(strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides),
		.agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality(strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality),
		.agg_sram_shared_loops_in2buf_autovec_write_0_ranges(strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges),
		.agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality(strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality),
		.agg_sram_shared_loops_in2buf_autovec_write_1_ranges(strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges),
		.chain_chain_en(strg_ub_vec_inst_chain_chain_en),
		.chain_data_in(strg_ub_vec_inst_chain_data_in),
		.clk(clk),
		.clk_en(clk_en),
		.data_from_strg(data_from_strg_lifted),
		.data_in(strg_ub_vec_inst_data_in),
		.flush(flush),
		.rst_n(rst_n),
		.sram_only_input_addr_gen_0_starting_addr(strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr),
		.sram_only_input_addr_gen_0_strides(strg_ub_vec_inst_sram_only_input_addr_gen_0_strides),
		.sram_only_input_addr_gen_1_starting_addr(strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr),
		.sram_only_input_addr_gen_1_strides(strg_ub_vec_inst_sram_only_input_addr_gen_1_strides),
		.sram_only_output_addr_gen_0_starting_addr(strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr),
		.sram_only_output_addr_gen_0_strides(strg_ub_vec_inst_sram_only_output_addr_gen_0_strides),
		.sram_only_output_addr_gen_1_starting_addr(strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr),
		.sram_only_output_addr_gen_1_strides(strg_ub_vec_inst_sram_only_output_addr_gen_1_strides),
		// .sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality),
		// .sram_tb_shared_loops_buf2out_autovec_read_0_ranges(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges),
		// .sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality),
		// .sram_tb_shared_loops_buf2out_autovec_read_1_ranges(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges),
		// .sram_tb_shared_output_sched_gen_0_enable(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable),
		// .sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr),
		// .sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides),
		// .sram_tb_shared_output_sched_gen_1_enable(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable),
		// .sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr),
		// .sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides),
		// .tb_only_loops_buf2out_read_0_dimensionality(strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality),
		// .tb_only_loops_buf2out_read_0_ranges(strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges),
		// .tb_only_loops_buf2out_read_1_dimensionality(strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality),
		// .tb_only_loops_buf2out_read_1_ranges(strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges),
		// .tb_only_tb_read_addr_gen_0_starting_addr(strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr),
		// .tb_only_tb_read_addr_gen_0_strides(strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides),
		// .tb_only_tb_read_addr_gen_1_starting_addr(strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr),
		// .tb_only_tb_read_addr_gen_1_strides(strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides),
		// .tb_only_tb_read_sched_gen_0_enable(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable),
		// .tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr),
		// .tb_only_tb_read_sched_gen_0_sched_addr_gen_strides(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides),
		// .tb_only_tb_read_sched_gen_1_enable(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable),
		// .tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr),
		// .tb_only_tb_read_sched_gen_1_sched_addr_gen_strides(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides),
		// .tb_only_tb_write_addr_gen_0_starting_addr(strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr),
		// .tb_only_tb_write_addr_gen_0_strides(strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides),
		// .tb_only_tb_write_addr_gen_1_starting_addr(strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr),
		// .tb_only_tb_write_addr_gen_1_strides(strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides),
		.accessor_output(strg_ub_vec_inst_accessor_output),
		.data_out(strg_ub_vec_inst_data_out),
		.data_to_strg(data_to_strg_lifted),
		.rd_addr_out(rd_addr_out_lifted),
		.ren_to_strg(ren_to_strg_lifted),
		.tmp0_rdaddr(tmp0_rdaddr_lifted),
		.tmp0_rden(tmp0_rden_lifted),
		.wen_to_strg(wen_to_strg_lifted),
		.wr_addr_out(wr_addr_out_lifted)
	);
endmodule
module LUT (
	lut,
	bit0,
	bit1,
	bit2,
	O,
	CLK,
	ASYNCRESET
);
	input [7:0] lut;
	input bit0;
	input bit1;
	input bit2;
	output O;
	input CLK;
	input ASYNCRESET;
	wire bit_const_0_None_out;
	wire [7:0] const_1_8_out;
	wire [7:0] magma_Bits_8_and_inst0_out;
	wire [7:0] magma_Bits_8_lshr_inst0_out;
	corebit_const #(.value(1'b0)) bit_const_0_None(.out(bit_const_0_None_out));
	coreir_const #(
		.value(8'h01),
		.width(8)
	) const_1_8(.out(const_1_8_out));
	coreir_and #(.width(8)) magma_Bits_8_and_inst0(
		.in0(magma_Bits_8_lshr_inst0_out),
		.in1(const_1_8_out),
		.out(magma_Bits_8_and_inst0_out)
	);
	wire [7:0] magma_Bits_8_lshr_inst0_in1;
	assign magma_Bits_8_lshr_inst0_in1 = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit2, bit1, bit0};
	coreir_lshr #(.width(8)) magma_Bits_8_lshr_inst0(
		.in0(lut),
		.in1(magma_Bits_8_lshr_inst0_in1),
		.out(magma_Bits_8_lshr_inst0_out)
	);
	assign O = magma_Bits_8_and_inst0_out[0];
endmodule
module Decode98 (
	I,
	O
);
	input [7:0] I;
	output O;
	wire [7:0] const_9_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h09),
		.width(8)
	) const_9_8(.out(const_9_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_9_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode88 (
	I,
	O
);
	input [7:0] I;
	output O;
	wire [7:0] const_8_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h08),
		.width(8)
	) const_8_8(.out(const_8_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_8_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode78 (
	I,
	O
);
	input [7:0] I;
	output O;
	wire [7:0] const_7_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h07),
		.width(8)
	) const_7_8(.out(const_7_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_7_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode68 (
	I,
	O
);
	input [7:0] I;
	output O;
	wire [7:0] const_6_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h06),
		.width(8)
	) const_6_8(.out(const_6_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_6_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode58 (
	I,
	O
);
	input [7:0] I;
	output O;
	wire [7:0] const_5_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h05),
		.width(8)
	) const_5_8(.out(const_5_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_5_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode48 (
	I,
	O
);
	input [7:0] I;
	output O;
	wire [7:0] const_4_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h04),
		.width(8)
	) const_4_8(.out(const_4_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_4_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode38 (
	I,
	O
);
	input [7:0] I;
	output O;
	wire [7:0] const_3_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h03),
		.width(8)
	) const_3_8(.out(const_3_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_3_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode28 (
	I,
	O
);
	input [7:0] I;
	output O;
	wire [7:0] const_2_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h02),
		.width(8)
	) const_2_8(.out(const_2_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_2_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode18 (
	I,
	O
);
	input [7:0] I;
	output O;
	wire [7:0] const_1_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h01),
		.width(8)
	) const_1_8(.out(const_1_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_1_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode108 (
	I,
	O
);
	input [7:0] I;
	output O;
	wire [7:0] const_10_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h0a),
		.width(8)
	) const_10_8(.out(const_10_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_10_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module Decode08 (
	I,
	O
);
	input [7:0] I;
	output O;
	wire [7:0] const_0_8_out;
	wire coreir_eq_8_inst0_out;
	coreir_const #(
		.value(8'h00),
		.width(8)
	) const_0_8(.out(const_0_8_out));
	coreir_eq #(.width(8)) coreir_eq_8_inst0(
		.in0(I),
		.in1(const_0_8_out),
		.out(coreir_eq_8_inst0_out)
	);
	assign O = coreir_eq_8_inst0_out;
endmodule
module ConfigRegister_4_8_32_1 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [3:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [3:0] Register_inst0_O;
	wire [7:0] const_1_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data[3:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h01),
		.width(8)
	) const_1_8(.out(const_1_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_1_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_4_8_32_0 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [3:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [3:0] Register_inst0_O;
	wire [7:0] const_0_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register Register_inst0(
		.I(config_data[3:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h00),
		.width(8)
	) const_0_8(.out(const_0_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_0_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_9 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_9_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h09),
		.width(8)
	) const_9_8(.out(const_9_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_9_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_80 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_80_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h50),
		.width(8)
	) const_80_8(.out(const_80_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_80_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_8 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_8_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h08),
		.width(8)
	) const_8_8(.out(const_8_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_8_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_79 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_79_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h4f),
		.width(8)
	) const_79_8(.out(const_79_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_79_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_78 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_78_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h4e),
		.width(8)
	) const_78_8(.out(const_78_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_78_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_77 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_77_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h4d),
		.width(8)
	) const_77_8(.out(const_77_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_77_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_76 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_76_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h4c),
		.width(8)
	) const_76_8(.out(const_76_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_76_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_74 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_74_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h4a),
		.width(8)
	) const_74_8(.out(const_74_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_74_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_73 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_73_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h49),
		.width(8)
	) const_73_8(.out(const_73_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_73_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_72 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_72_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h48),
		.width(8)
	) const_72_8(.out(const_72_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_72_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_70 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_70_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h46),
		.width(8)
	) const_70_8(.out(const_70_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_70_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_7 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_7_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h07),
		.width(8)
	) const_7_8(.out(const_7_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_7_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_69 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_69_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h45),
		.width(8)
	) const_69_8(.out(const_69_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_69_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_68 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_68_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h44),
		.width(8)
	) const_68_8(.out(const_68_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_68_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_67 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_67_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h43),
		.width(8)
	) const_67_8(.out(const_67_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_67_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_65 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_65_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h41),
		.width(8)
	) const_65_8(.out(const_65_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_65_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_64 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_64_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h40),
		.width(8)
	) const_64_8(.out(const_64_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_64_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_62 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_62_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h3e),
		.width(8)
	) const_62_8(.out(const_62_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_62_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_61 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_61_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h3d),
		.width(8)
	) const_61_8(.out(const_61_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_61_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_60 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_60_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h3c),
		.width(8)
	) const_60_8(.out(const_60_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_60_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_6 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_6_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h06),
		.width(8)
	) const_6_8(.out(const_6_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_6_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_58 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_58_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h3a),
		.width(8)
	) const_58_8(.out(const_58_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_58_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_57 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_57_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h39),
		.width(8)
	) const_57_8(.out(const_57_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_57_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_56 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_56_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h38),
		.width(8)
	) const_56_8(.out(const_56_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_56_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_54 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_54_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h36),
		.width(8)
	) const_54_8(.out(const_54_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_54_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_53 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_53_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h35),
		.width(8)
	) const_53_8(.out(const_53_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_53_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_52 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_52_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h34),
		.width(8)
	) const_52_8(.out(const_52_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_52_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_50 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_50_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h32),
		.width(8)
	) const_50_8(.out(const_50_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_50_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_5 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_5_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h05),
		.width(8)
	) const_5_8(.out(const_5_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_5_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_49 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_49_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h31),
		.width(8)
	) const_49_8(.out(const_49_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_49_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_47 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_47_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h2f),
		.width(8)
	) const_47_8(.out(const_47_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_47_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_46 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_46_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h2e),
		.width(8)
	) const_46_8(.out(const_46_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_46_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_45 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_45_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h2d),
		.width(8)
	) const_45_8(.out(const_45_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_45_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_44 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_44_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h2c),
		.width(8)
	) const_44_8(.out(const_44_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_44_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_43 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_43_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h2b),
		.width(8)
	) const_43_8(.out(const_43_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_43_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_42 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_42_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h2a),
		.width(8)
	) const_42_8(.out(const_42_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_42_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_40 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_40_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h28),
		.width(8)
	) const_40_8(.out(const_40_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_40_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_4 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_4_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h04),
		.width(8)
	) const_4_8(.out(const_4_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_4_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_39 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_39_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h27),
		.width(8)
	) const_39_8(.out(const_39_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_39_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_38 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_38_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h26),
		.width(8)
	) const_38_8(.out(const_38_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_38_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_36 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_36_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h24),
		.width(8)
	) const_36_8(.out(const_36_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_36_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_35 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_35_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h23),
		.width(8)
	) const_35_8(.out(const_35_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_35_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_33 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_33_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h21),
		.width(8)
	) const_33_8(.out(const_33_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_33_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_32 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_32_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h20),
		.width(8)
	) const_32_8(.out(const_32_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_32_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_31 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_31_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h1f),
		.width(8)
	) const_31_8(.out(const_31_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_31_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_29 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_29_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h1d),
		.width(8)
	) const_29_8(.out(const_29_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_29_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_28 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_28_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h1c),
		.width(8)
	) const_28_8(.out(const_28_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_28_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_27 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_27_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h1b),
		.width(8)
	) const_27_8(.out(const_27_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_27_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_25 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_25_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h19),
		.width(8)
	) const_25_8(.out(const_25_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_25_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_24 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_24_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h18),
		.width(8)
	) const_24_8(.out(const_24_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_24_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_23 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_23_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h17),
		.width(8)
	) const_23_8(.out(const_23_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_23_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_21 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_21_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h15),
		.width(8)
	) const_21_8(.out(const_21_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_21_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_20 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_20_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h14),
		.width(8)
	) const_20_8(.out(const_20_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_20_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_2 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_2_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h02),
		.width(8)
	) const_2_8(.out(const_2_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_2_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_18 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_18_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h12),
		.width(8)
	) const_18_8(.out(const_18_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_18_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_17 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_17_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h11),
		.width(8)
	) const_17_8(.out(const_17_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_17_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_16 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_16_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h10),
		.width(8)
	) const_16_8(.out(const_16_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_16_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_14 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_14_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h0e),
		.width(8)
	) const_14_8(.out(const_14_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_14_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_13 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_13_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h0d),
		.width(8)
	) const_13_8(.out(const_13_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_13_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_12 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_12_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h0c),
		.width(8)
	) const_12_8(.out(const_12_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_12_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_10 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_10_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h0a),
		.width(8)
	) const_10_8(.out(const_10_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_10_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_1 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_1_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h01),
		.width(8)
	) const_1_8(.out(const_1_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_1_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_32_8_32_0 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [31:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [31:0] Register_inst0_O;
	wire [7:0] const_0_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq3 Register_inst0(
		.I(config_data),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h00),
		.width(8)
	) const_0_8(.out(const_0_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_0_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module SB_ID0_3TRACKS_B1_PE (
	SB_T0_EAST_SB_IN_B1,
	SB_T0_EAST_SB_OUT_B1,
	SB_T0_NORTH_SB_IN_B1,
	SB_T0_NORTH_SB_OUT_B1,
	SB_T0_SOUTH_SB_IN_B1,
	SB_T0_SOUTH_SB_OUT_B1,
	SB_T0_WEST_SB_IN_B1,
	SB_T0_WEST_SB_OUT_B1,
	SB_T1_EAST_SB_IN_B1,
	SB_T1_EAST_SB_OUT_B1,
	SB_T1_NORTH_SB_IN_B1,
	SB_T1_NORTH_SB_OUT_B1,
	SB_T1_SOUTH_SB_IN_B1,
	SB_T1_SOUTH_SB_OUT_B1,
	SB_T1_WEST_SB_IN_B1,
	SB_T1_WEST_SB_OUT_B1,
	SB_T2_EAST_SB_IN_B1,
	SB_T2_EAST_SB_OUT_B1,
	SB_T2_NORTH_SB_IN_B1,
	SB_T2_NORTH_SB_OUT_B1,
	SB_T2_SOUTH_SB_IN_B1,
	SB_T2_SOUTH_SB_OUT_B1,
	SB_T2_WEST_SB_IN_B1,
	SB_T2_WEST_SB_OUT_B1,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	read_config_data,
	res_p,
	reset,
	stall
);
	input [0:0] SB_T0_EAST_SB_IN_B1;
	output [0:0] SB_T0_EAST_SB_OUT_B1;
	input [0:0] SB_T0_NORTH_SB_IN_B1;
	output [0:0] SB_T0_NORTH_SB_OUT_B1;
	input [0:0] SB_T0_SOUTH_SB_IN_B1;
	output [0:0] SB_T0_SOUTH_SB_OUT_B1;
	input [0:0] SB_T0_WEST_SB_IN_B1;
	output [0:0] SB_T0_WEST_SB_OUT_B1;
	input [0:0] SB_T1_EAST_SB_IN_B1;
	output [0:0] SB_T1_EAST_SB_OUT_B1;
	input [0:0] SB_T1_NORTH_SB_IN_B1;
	output [0:0] SB_T1_NORTH_SB_OUT_B1;
	input [0:0] SB_T1_SOUTH_SB_IN_B1;
	output [0:0] SB_T1_SOUTH_SB_OUT_B1;
	input [0:0] SB_T1_WEST_SB_IN_B1;
	output [0:0] SB_T1_WEST_SB_OUT_B1;
	input [0:0] SB_T2_EAST_SB_IN_B1;
	output [0:0] SB_T2_EAST_SB_OUT_B1;
	input [0:0] SB_T2_NORTH_SB_IN_B1;
	output [0:0] SB_T2_NORTH_SB_OUT_B1;
	input [0:0] SB_T2_SOUTH_SB_IN_B1;
	output [0:0] SB_T2_SOUTH_SB_OUT_B1;
	input [0:0] SB_T2_WEST_SB_IN_B1;
	output [0:0] SB_T2_WEST_SB_OUT_B1;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output [31:0] read_config_data;
	input [0:0] res_p;
	input reset;
	input [0:0] stall;
	wire [0:0] Invert1_inst0_out;
	wire [0:0] MUX_SB_T0_EAST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out;
	wire [0:0] MUX_SB_T0_NORTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out;
	wire [0:0] MUX_SB_T0_SOUTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out;
	wire [0:0] MUX_SB_T0_WEST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out;
	wire [0:0] MUX_SB_T1_EAST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out;
	wire [0:0] MUX_SB_T1_NORTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out;
	wire [0:0] MUX_SB_T1_SOUTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out;
	wire [0:0] MUX_SB_T1_WEST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out;
	wire [0:0] MUX_SB_T2_EAST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out;
	wire [0:0] MUX_SB_T2_NORTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out;
	wire [0:0] MUX_SB_T2_SOUTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out;
	wire [0:0] MUX_SB_T2_WEST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out;
	wire [31:0] MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
	wire [0:0] REG_T0_EAST_B1_O;
	wire [0:0] REG_T0_NORTH_B1_O;
	wire [0:0] REG_T0_SOUTH_B1_O;
	wire [0:0] REG_T0_WEST_B1_O;
	wire [0:0] REG_T1_EAST_B1_O;
	wire [0:0] REG_T1_NORTH_B1_O;
	wire [0:0] REG_T1_SOUTH_B1_O;
	wire [0:0] REG_T1_WEST_B1_O;
	wire [0:0] REG_T2_EAST_B1_O;
	wire [0:0] REG_T2_NORTH_B1_O;
	wire [0:0] REG_T2_SOUTH_B1_O;
	wire [0:0] REG_T2_WEST_B1_O;
	wire [0:0] RMUX_T0_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T0_EAST_B1_sel_inst0_O;
	wire [0:0] RMUX_T0_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T0_NORTH_B1_sel_inst0_O;
	wire [0:0] RMUX_T0_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T0_SOUTH_B1_sel_inst0_O;
	wire [0:0] RMUX_T0_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T0_WEST_B1_sel_inst0_O;
	wire [0:0] RMUX_T1_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T1_EAST_B1_sel_inst0_O;
	wire [0:0] RMUX_T1_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T1_NORTH_B1_sel_inst0_O;
	wire [0:0] RMUX_T1_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T1_SOUTH_B1_sel_inst0_O;
	wire [0:0] RMUX_T1_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T1_WEST_B1_sel_inst0_O;
	wire [0:0] RMUX_T2_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T2_EAST_B1_sel_inst0_O;
	wire [0:0] RMUX_T2_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T2_NORTH_B1_sel_inst0_O;
	wire [0:0] RMUX_T2_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T2_SOUTH_B1_sel_inst0_O;
	wire [0:0] RMUX_T2_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T2_WEST_B1_sel_inst0_O;
	wire [1:0] SB_T0_EAST_SB_OUT_B1_sel_inst0_O;
	wire [1:0] SB_T0_NORTH_SB_OUT_B1_sel_inst0_O;
	wire [1:0] SB_T0_SOUTH_SB_OUT_B1_sel_inst0_O;
	wire [1:0] SB_T0_WEST_SB_OUT_B1_sel_inst0_O;
	wire [1:0] SB_T1_EAST_SB_OUT_B1_sel_inst0_O;
	wire [1:0] SB_T1_NORTH_SB_OUT_B1_sel_inst0_O;
	wire [1:0] SB_T1_SOUTH_SB_OUT_B1_sel_inst0_O;
	wire [1:0] SB_T1_WEST_SB_OUT_B1_sel_inst0_O;
	wire [1:0] SB_T2_EAST_SB_OUT_B1_sel_inst0_O;
	wire [1:0] SB_T2_NORTH_SB_OUT_B1_sel_inst0_O;
	wire [1:0] SB_T2_SOUTH_SB_OUT_B1_sel_inst0_O;
	wire [1:0] SB_T2_WEST_SB_OUT_B1_sel_inst0_O;
	wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1_O;
	wire ZextWrapper_4_32_inst0$bit_const_0_None_out;
	wire [3:0] ZextWrapper_4_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_4_32_inst0$self_O_in;
	wire [0:0] and1_inst0_out;
	wire [0:0] and1_inst1_out;
	wire [0:0] and1_inst10_out;
	wire [0:0] and1_inst11_out;
	wire [0:0] and1_inst2_out;
	wire [0:0] and1_inst3_out;
	wire [0:0] and1_inst4_out;
	wire [0:0] and1_inst5_out;
	wire [0:0] and1_inst6_out;
	wire [0:0] and1_inst7_out;
	wire [0:0] and1_inst8_out;
	wire [0:0] and1_inst9_out;
	wire [31:0] config_reg_0_O;
	wire [3:0] config_reg_1_O;
	wire [0:0] const_1_1_out;
	wire coreir_eq_1_inst0_out;
	wire coreir_eq_1_inst1_out;
	wire coreir_eq_1_inst10_out;
	wire coreir_eq_1_inst11_out;
	wire coreir_eq_1_inst2_out;
	wire coreir_eq_1_inst3_out;
	wire coreir_eq_1_inst4_out;
	wire coreir_eq_1_inst5_out;
	wire coreir_eq_1_inst6_out;
	wire coreir_eq_1_inst7_out;
	wire coreir_eq_1_inst8_out;
	wire coreir_eq_1_inst9_out;
	coreir_not #(.width(1)) Invert1_inst0(
		.in(stall),
		.out(Invert1_inst0_out)
	);
	commonlib_muxn__N4__width1 MUX_SB_T0_EAST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0(
		.in_data_0(WIRE_SB_T0_WEST_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T2_NORTH_SB_IN_B1_O),
		.in_data_3(res_p),
		.in_sel(SB_T0_EAST_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T0_EAST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out)
	);
	commonlib_muxn__N4__width1 MUX_SB_T0_NORTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0(
		.in_data_0(WIRE_SB_T0_WEST_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T1_EAST_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
		.in_data_3(res_p),
		.in_sel(SB_T0_NORTH_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T0_NORTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out)
	);
	commonlib_muxn__N4__width1 MUX_SB_T0_SOUTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0(
		.in_data_0(WIRE_SB_T1_EAST_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T0_NORTH_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T1_WEST_SB_IN_B1_O),
		.in_data_3(res_p),
		.in_sel(SB_T0_SOUTH_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T0_SOUTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out)
	);
	commonlib_muxn__N4__width1 MUX_SB_T0_WEST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0(
		.in_data_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
		.in_data_3(res_p),
		.in_sel(SB_T0_WEST_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T0_WEST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out)
	);
	commonlib_muxn__N4__width1 MUX_SB_T1_EAST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0(
		.in_data_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T1_WEST_SB_IN_B1_O),
		.in_data_3(res_p),
		.in_sel(SB_T1_EAST_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T1_EAST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out)
	);
	commonlib_muxn__N4__width1 MUX_SB_T1_NORTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0(
		.in_data_0(WIRE_SB_T2_EAST_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T2_WEST_SB_IN_B1_O),
		.in_data_3(res_p),
		.in_sel(SB_T1_NORTH_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T1_NORTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out)
	);
	commonlib_muxn__N4__width1 MUX_SB_T1_SOUTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0(
		.in_data_0(WIRE_SB_T0_EAST_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T1_NORTH_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T2_WEST_SB_IN_B1_O),
		.in_data_3(res_p),
		.in_sel(SB_T1_SOUTH_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T1_SOUTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out)
	);
	commonlib_muxn__N4__width1 MUX_SB_T1_WEST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0(
		.in_data_0(WIRE_SB_T2_NORTH_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T1_EAST_SB_IN_B1_O),
		.in_data_3(res_p),
		.in_sel(SB_T1_WEST_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T1_WEST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out)
	);
	commonlib_muxn__N4__width1 MUX_SB_T2_EAST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0(
		.in_data_0(WIRE_SB_T1_NORTH_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T2_WEST_SB_IN_B1_O),
		.in_data_3(res_p),
		.in_sel(SB_T2_EAST_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T2_EAST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out)
	);
	commonlib_muxn__N4__width1 MUX_SB_T2_NORTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0(
		.in_data_0(WIRE_SB_T1_WEST_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T0_EAST_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
		.in_data_3(res_p),
		.in_sel(SB_T2_NORTH_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T2_NORTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out)
	);
	commonlib_muxn__N4__width1 MUX_SB_T2_SOUTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0(
		.in_data_0(WIRE_SB_T0_WEST_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T2_EAST_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T2_NORTH_SB_IN_B1_O),
		.in_data_3(res_p),
		.in_sel(SB_T2_SOUTH_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T2_SOUTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out)
	);
	commonlib_muxn__N4__width1 MUX_SB_T2_WEST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0(
		.in_data_0(WIRE_SB_T1_NORTH_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T2_EAST_SB_IN_B1_O),
		.in_data_3(res_p),
		.in_sel(SB_T2_WEST_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T2_WEST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out)
	);
	coreir_mux #(.width(32)) MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join(
		.in0(config_reg_0_O),
		.in1(ZextWrapper_4_32_inst0$self_O_in),
		.sel(config_config_addr[0]),
		.out(MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out)
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_EAST_B1(
		.I(MUX_SB_T0_EAST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.O(REG_T0_EAST_B1_O),
		.CLK(clk),
		.CE(and1_inst2_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_NORTH_B1(
		.I(MUX_SB_T0_NORTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.O(REG_T0_NORTH_B1_O),
		.CLK(clk),
		.CE(and1_inst0_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_SOUTH_B1(
		.I(MUX_SB_T0_SOUTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.O(REG_T0_SOUTH_B1_O),
		.CLK(clk),
		.CE(and1_inst1_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_WEST_B1(
		.I(MUX_SB_T0_WEST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.O(REG_T0_WEST_B1_O),
		.CLK(clk),
		.CE(and1_inst3_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_EAST_B1(
		.I(MUX_SB_T1_EAST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.O(REG_T1_EAST_B1_O),
		.CLK(clk),
		.CE(and1_inst6_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_NORTH_B1(
		.I(MUX_SB_T1_NORTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.O(REG_T1_NORTH_B1_O),
		.CLK(clk),
		.CE(and1_inst4_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_SOUTH_B1(
		.I(MUX_SB_T1_SOUTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.O(REG_T1_SOUTH_B1_O),
		.CLK(clk),
		.CE(and1_inst5_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_WEST_B1(
		.I(MUX_SB_T1_WEST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.O(REG_T1_WEST_B1_O),
		.CLK(clk),
		.CE(and1_inst7_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_EAST_B1(
		.I(MUX_SB_T2_EAST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.O(REG_T2_EAST_B1_O),
		.CLK(clk),
		.CE(and1_inst10_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_NORTH_B1(
		.I(MUX_SB_T2_NORTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.O(REG_T2_NORTH_B1_O),
		.CLK(clk),
		.CE(and1_inst8_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_SOUTH_B1(
		.I(MUX_SB_T2_SOUTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.O(REG_T2_SOUTH_B1_O),
		.CLK(clk),
		.CE(and1_inst9_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_WEST_B1(
		.I(MUX_SB_T2_WEST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.O(REG_T2_WEST_B1_O),
		.CLK(clk),
		.CE(and1_inst11_out[0])
	);
	coreir_mux #(.width(1)) RMUX_T0_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T0_EAST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.in1(REG_T0_EAST_B1_O),
		.sel(RMUX_T0_EAST_B1_sel_inst0_O[0]),
		.out(RMUX_T0_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T0_EAST_B1_sel RMUX_T0_EAST_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T0_EAST_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T0_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T0_NORTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.in1(REG_T0_NORTH_B1_O),
		.sel(RMUX_T0_NORTH_B1_sel_inst0_O[0]),
		.out(RMUX_T0_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T0_NORTH_B1_sel RMUX_T0_NORTH_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T0_NORTH_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T0_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T0_SOUTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.in1(REG_T0_SOUTH_B1_O),
		.sel(RMUX_T0_SOUTH_B1_sel_inst0_O[0]),
		.out(RMUX_T0_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T0_SOUTH_B1_sel RMUX_T0_SOUTH_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T0_SOUTH_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T0_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T0_WEST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.in1(REG_T0_WEST_B1_O),
		.sel(RMUX_T0_WEST_B1_sel_inst0_O[0]),
		.out(RMUX_T0_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T0_WEST_B1_sel RMUX_T0_WEST_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T0_WEST_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T1_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T1_EAST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.in1(REG_T1_EAST_B1_O),
		.sel(RMUX_T1_EAST_B1_sel_inst0_O[0]),
		.out(RMUX_T1_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T1_EAST_B1_sel RMUX_T1_EAST_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T1_EAST_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T1_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T1_NORTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.in1(REG_T1_NORTH_B1_O),
		.sel(RMUX_T1_NORTH_B1_sel_inst0_O[0]),
		.out(RMUX_T1_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T1_NORTH_B1_sel RMUX_T1_NORTH_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T1_NORTH_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T1_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T1_SOUTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.in1(REG_T1_SOUTH_B1_O),
		.sel(RMUX_T1_SOUTH_B1_sel_inst0_O[0]),
		.out(RMUX_T1_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T1_SOUTH_B1_sel RMUX_T1_SOUTH_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T1_SOUTH_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T1_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T1_WEST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.in1(REG_T1_WEST_B1_O),
		.sel(RMUX_T1_WEST_B1_sel_inst0_O[0]),
		.out(RMUX_T1_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T1_WEST_B1_sel RMUX_T1_WEST_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T1_WEST_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T2_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T2_EAST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.in1(REG_T2_EAST_B1_O),
		.sel(RMUX_T2_EAST_B1_sel_inst0_O[0]),
		.out(RMUX_T2_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T2_EAST_B1_sel RMUX_T2_EAST_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T2_EAST_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T2_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T2_NORTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.in1(REG_T2_NORTH_B1_O),
		.sel(RMUX_T2_NORTH_B1_sel_inst0_O[0]),
		.out(RMUX_T2_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T2_NORTH_B1_sel RMUX_T2_NORTH_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T2_NORTH_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T2_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T2_SOUTH_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.in1(REG_T2_SOUTH_B1_O),
		.sel(RMUX_T2_SOUTH_B1_sel_inst0_O[0]),
		.out(RMUX_T2_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T2_SOUTH_B1_sel RMUX_T2_SOUTH_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T2_SOUTH_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T2_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T2_WEST_SB_OUT_B1$Mux4xBits1_inst0$coreir_commonlib_mux4x1_inst0_out),
		.in1(REG_T2_WEST_B1_O),
		.sel(RMUX_T2_WEST_B1_sel_inst0_O[0]),
		.out(RMUX_T2_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T2_WEST_B1_sel RMUX_T2_WEST_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T2_WEST_B1_sel_inst0_O)
	);
	SB_T0_EAST_SB_OUT_B1_sel SB_T0_EAST_SB_OUT_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T0_EAST_SB_OUT_B1_sel_inst0_O)
	);
	SB_T0_NORTH_SB_OUT_B1_sel SB_T0_NORTH_SB_OUT_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T0_NORTH_SB_OUT_B1_sel_inst0_O)
	);
	SB_T0_SOUTH_SB_OUT_B1_sel SB_T0_SOUTH_SB_OUT_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T0_SOUTH_SB_OUT_B1_sel_inst0_O)
	);
	SB_T0_WEST_SB_OUT_B1_sel SB_T0_WEST_SB_OUT_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T0_WEST_SB_OUT_B1_sel_inst0_O)
	);
	SB_T1_EAST_SB_OUT_B1_sel SB_T1_EAST_SB_OUT_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T1_EAST_SB_OUT_B1_sel_inst0_O)
	);
	SB_T1_NORTH_SB_OUT_B1_sel SB_T1_NORTH_SB_OUT_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T1_NORTH_SB_OUT_B1_sel_inst0_O)
	);
	SB_T1_SOUTH_SB_OUT_B1_sel SB_T1_SOUTH_SB_OUT_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T1_SOUTH_SB_OUT_B1_sel_inst0_O)
	);
	SB_T1_WEST_SB_OUT_B1_sel SB_T1_WEST_SB_OUT_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T1_WEST_SB_OUT_B1_sel_inst0_O)
	);
	SB_T2_EAST_SB_OUT_B1_sel SB_T2_EAST_SB_OUT_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T2_EAST_SB_OUT_B1_sel_inst0_O)
	);
	SB_T2_NORTH_SB_OUT_B1_sel SB_T2_NORTH_SB_OUT_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T2_NORTH_SB_OUT_B1_sel_inst0_O)
	);
	SB_T2_SOUTH_SB_OUT_B1_sel SB_T2_SOUTH_SB_OUT_B1_sel_inst0(
		.I(config_reg_1_O),
		.O(SB_T2_SOUTH_SB_OUT_B1_sel_inst0_O)
	);
	SB_T2_WEST_SB_OUT_B1_sel SB_T2_WEST_SB_OUT_B1_sel_inst0(
		.I(config_reg_1_O),
		.O(SB_T2_WEST_SB_OUT_B1_sel_inst0_O)
	);
	MuxWrapper_1_1 WIRE_SB_T0_EAST_SB_IN_B1(
		.I(SB_T0_EAST_SB_IN_B1),
		.O(WIRE_SB_T0_EAST_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T0_NORTH_SB_IN_B1(
		.I(SB_T0_NORTH_SB_IN_B1),
		.O(WIRE_SB_T0_NORTH_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T0_SOUTH_SB_IN_B1(
		.I(SB_T0_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T0_SOUTH_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T0_WEST_SB_IN_B1(
		.I(SB_T0_WEST_SB_IN_B1),
		.O(WIRE_SB_T0_WEST_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T1_EAST_SB_IN_B1(
		.I(SB_T1_EAST_SB_IN_B1),
		.O(WIRE_SB_T1_EAST_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T1_NORTH_SB_IN_B1(
		.I(SB_T1_NORTH_SB_IN_B1),
		.O(WIRE_SB_T1_NORTH_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T1_SOUTH_SB_IN_B1(
		.I(SB_T1_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T1_SOUTH_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T1_WEST_SB_IN_B1(
		.I(SB_T1_WEST_SB_IN_B1),
		.O(WIRE_SB_T1_WEST_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T2_EAST_SB_IN_B1(
		.I(SB_T2_EAST_SB_IN_B1),
		.O(WIRE_SB_T2_EAST_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T2_NORTH_SB_IN_B1(
		.I(SB_T2_NORTH_SB_IN_B1),
		.O(WIRE_SB_T2_NORTH_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T2_SOUTH_SB_IN_B1(
		.I(SB_T2_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T2_SOUTH_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T2_WEST_SB_IN_B1(
		.I(SB_T2_WEST_SB_IN_B1),
		.O(WIRE_SB_T2_WEST_SB_IN_B1_O)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_4_32_inst0$bit_const_0_None(.out(ZextWrapper_4_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit4 ZextWrapper_4_32_inst0$self_I(
		.in(config_reg_1_O),
		.out(ZextWrapper_4_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_4_32_inst0$self_O_out;
	assign ZextWrapper_4_32_inst0$self_O_out = {ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$self_I_out[3:0]};
	mantle_wire__typeBitIn32 ZextWrapper_4_32_inst0$self_O(
		.in(ZextWrapper_4_32_inst0$self_O_in),
		.out(ZextWrapper_4_32_inst0$self_O_out)
	);
	coreir_and #(.width(1)) and1_inst0(
		.in0(coreir_eq_1_inst0_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst0_out)
	);
	coreir_and #(.width(1)) and1_inst1(
		.in0(coreir_eq_1_inst1_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst1_out)
	);
	coreir_and #(.width(1)) and1_inst10(
		.in0(coreir_eq_1_inst10_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst10_out)
	);
	coreir_and #(.width(1)) and1_inst11(
		.in0(coreir_eq_1_inst11_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst11_out)
	);
	coreir_and #(.width(1)) and1_inst2(
		.in0(coreir_eq_1_inst2_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst2_out)
	);
	coreir_and #(.width(1)) and1_inst3(
		.in0(coreir_eq_1_inst3_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst3_out)
	);
	coreir_and #(.width(1)) and1_inst4(
		.in0(coreir_eq_1_inst4_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst4_out)
	);
	coreir_and #(.width(1)) and1_inst5(
		.in0(coreir_eq_1_inst5_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst5_out)
	);
	coreir_and #(.width(1)) and1_inst6(
		.in0(coreir_eq_1_inst6_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst6_out)
	);
	coreir_and #(.width(1)) and1_inst7(
		.in0(coreir_eq_1_inst7_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst7_out)
	);
	coreir_and #(.width(1)) and1_inst8(
		.in0(coreir_eq_1_inst8_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst8_out)
	);
	coreir_and #(.width(1)) and1_inst9(
		.in0(coreir_eq_1_inst9_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst9_out)
	);
	ConfigRegister_32_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_4_8_32_1 config_reg_1(
		.clk(clk),
		.reset(reset),
		.O(config_reg_1_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	coreir_const #(
		.value(1'h1),
		.width(1)
	) const_1_1(.out(const_1_1_out));
	coreir_eq #(.width(1)) coreir_eq_1_inst0(
		.in0(const_1_1_out),
		.in1(RMUX_T0_NORTH_B1_sel_inst0_O),
		.out(coreir_eq_1_inst0_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst1(
		.in0(const_1_1_out),
		.in1(RMUX_T0_SOUTH_B1_sel_inst0_O),
		.out(coreir_eq_1_inst1_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst10(
		.in0(const_1_1_out),
		.in1(RMUX_T2_EAST_B1_sel_inst0_O),
		.out(coreir_eq_1_inst10_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst11(
		.in0(const_1_1_out),
		.in1(RMUX_T2_WEST_B1_sel_inst0_O),
		.out(coreir_eq_1_inst11_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst2(
		.in0(const_1_1_out),
		.in1(RMUX_T0_EAST_B1_sel_inst0_O),
		.out(coreir_eq_1_inst2_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst3(
		.in0(const_1_1_out),
		.in1(RMUX_T0_WEST_B1_sel_inst0_O),
		.out(coreir_eq_1_inst3_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst4(
		.in0(const_1_1_out),
		.in1(RMUX_T1_NORTH_B1_sel_inst0_O),
		.out(coreir_eq_1_inst4_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst5(
		.in0(const_1_1_out),
		.in1(RMUX_T1_SOUTH_B1_sel_inst0_O),
		.out(coreir_eq_1_inst5_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst6(
		.in0(const_1_1_out),
		.in1(RMUX_T1_EAST_B1_sel_inst0_O),
		.out(coreir_eq_1_inst6_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst7(
		.in0(const_1_1_out),
		.in1(RMUX_T1_WEST_B1_sel_inst0_O),
		.out(coreir_eq_1_inst7_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst8(
		.in0(const_1_1_out),
		.in1(RMUX_T2_NORTH_B1_sel_inst0_O),
		.out(coreir_eq_1_inst8_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst9(
		.in0(const_1_1_out),
		.in1(RMUX_T2_SOUTH_B1_sel_inst0_O),
		.out(coreir_eq_1_inst9_out)
	);
	assign SB_T0_EAST_SB_OUT_B1 = RMUX_T0_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T0_NORTH_SB_OUT_B1 = RMUX_T0_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T0_SOUTH_SB_OUT_B1 = RMUX_T0_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T0_WEST_SB_OUT_B1 = RMUX_T0_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T1_EAST_SB_OUT_B1 = RMUX_T1_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T1_NORTH_SB_OUT_B1 = RMUX_T1_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T1_SOUTH_SB_OUT_B1 = RMUX_T1_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T1_WEST_SB_OUT_B1 = RMUX_T1_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T2_EAST_SB_OUT_B1 = RMUX_T2_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T2_NORTH_SB_OUT_B1 = RMUX_T2_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T2_SOUTH_SB_OUT_B1 = RMUX_T2_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T2_WEST_SB_OUT_B1 = RMUX_T2_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign read_config_data = MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
endmodule
module SB_ID0_3TRACKS_B16_PE (
	SB_T0_EAST_SB_IN_B16,
	SB_T0_EAST_SB_OUT_B16,
	SB_T0_NORTH_SB_IN_B16,
	SB_T0_NORTH_SB_OUT_B16,
	SB_T0_SOUTH_SB_IN_B16,
	SB_T0_SOUTH_SB_OUT_B16,
	SB_T0_WEST_SB_IN_B16,
	SB_T0_WEST_SB_OUT_B16,
	SB_T1_EAST_SB_IN_B16,
	SB_T1_EAST_SB_OUT_B16,
	SB_T1_NORTH_SB_IN_B16,
	SB_T1_NORTH_SB_OUT_B16,
	SB_T1_SOUTH_SB_IN_B16,
	SB_T1_SOUTH_SB_OUT_B16,
	SB_T1_WEST_SB_IN_B16,
	SB_T1_WEST_SB_OUT_B16,
	SB_T2_EAST_SB_IN_B16,
	SB_T2_EAST_SB_OUT_B16,
	SB_T2_NORTH_SB_IN_B16,
	SB_T2_NORTH_SB_OUT_B16,
	SB_T2_SOUTH_SB_IN_B16,
	SB_T2_SOUTH_SB_OUT_B16,
	SB_T2_WEST_SB_IN_B16,
	SB_T2_WEST_SB_OUT_B16,
	alu_res,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	read_config_data,
	reset,
	stall
);
	input [15:0] SB_T0_EAST_SB_IN_B16;
	output [15:0] SB_T0_EAST_SB_OUT_B16;
	input [15:0] SB_T0_NORTH_SB_IN_B16;
	output [15:0] SB_T0_NORTH_SB_OUT_B16;
	input [15:0] SB_T0_SOUTH_SB_IN_B16;
	output [15:0] SB_T0_SOUTH_SB_OUT_B16;
	input [15:0] SB_T0_WEST_SB_IN_B16;
	output [15:0] SB_T0_WEST_SB_OUT_B16;
	input [15:0] SB_T1_EAST_SB_IN_B16;
	output [15:0] SB_T1_EAST_SB_OUT_B16;
	input [15:0] SB_T1_NORTH_SB_IN_B16;
	output [15:0] SB_T1_NORTH_SB_OUT_B16;
	input [15:0] SB_T1_SOUTH_SB_IN_B16;
	output [15:0] SB_T1_SOUTH_SB_OUT_B16;
	input [15:0] SB_T1_WEST_SB_IN_B16;
	output [15:0] SB_T1_WEST_SB_OUT_B16;
	input [15:0] SB_T2_EAST_SB_IN_B16;
	output [15:0] SB_T2_EAST_SB_OUT_B16;
	input [15:0] SB_T2_NORTH_SB_IN_B16;
	output [15:0] SB_T2_NORTH_SB_OUT_B16;
	input [15:0] SB_T2_SOUTH_SB_IN_B16;
	output [15:0] SB_T2_SOUTH_SB_OUT_B16;
	input [15:0] SB_T2_WEST_SB_IN_B16;
	output [15:0] SB_T2_WEST_SB_OUT_B16;
	input [15:0] alu_res;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output [31:0] read_config_data;
	input reset;
	input [0:0] stall;
	wire [0:0] Invert1_inst0_out;
	wire [15:0] MUX_SB_T0_EAST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out;
	wire [15:0] MUX_SB_T0_NORTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out;
	wire [15:0] MUX_SB_T0_SOUTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out;
	wire [15:0] MUX_SB_T0_WEST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out;
	wire [15:0] MUX_SB_T1_EAST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out;
	wire [15:0] MUX_SB_T1_NORTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out;
	wire [15:0] MUX_SB_T1_SOUTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out;
	wire [15:0] MUX_SB_T1_WEST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out;
	wire [15:0] MUX_SB_T2_EAST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out;
	wire [15:0] MUX_SB_T2_NORTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out;
	wire [15:0] MUX_SB_T2_SOUTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out;
	wire [15:0] MUX_SB_T2_WEST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out;
	wire [31:0] MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
	wire [15:0] REG_T0_EAST_B16_O;
	wire [15:0] REG_T0_NORTH_B16_O;
	wire [15:0] REG_T0_SOUTH_B16_O;
	wire [15:0] REG_T0_WEST_B16_O;
	wire [15:0] REG_T1_EAST_B16_O;
	wire [15:0] REG_T1_NORTH_B16_O;
	wire [15:0] REG_T1_SOUTH_B16_O;
	wire [15:0] REG_T1_WEST_B16_O;
	wire [15:0] REG_T2_EAST_B16_O;
	wire [15:0] REG_T2_NORTH_B16_O;
	wire [15:0] REG_T2_SOUTH_B16_O;
	wire [15:0] REG_T2_WEST_B16_O;
	wire [15:0] RMUX_T0_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T0_EAST_B16_sel_inst0_O;
	wire [15:0] RMUX_T0_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T0_NORTH_B16_sel_inst0_O;
	wire [15:0] RMUX_T0_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T0_SOUTH_B16_sel_inst0_O;
	wire [15:0] RMUX_T0_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T0_WEST_B16_sel_inst0_O;
	wire [15:0] RMUX_T1_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T1_EAST_B16_sel_inst0_O;
	wire [15:0] RMUX_T1_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T1_NORTH_B16_sel_inst0_O;
	wire [15:0] RMUX_T1_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T1_SOUTH_B16_sel_inst0_O;
	wire [15:0] RMUX_T1_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T1_WEST_B16_sel_inst0_O;
	wire [15:0] RMUX_T2_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T2_EAST_B16_sel_inst0_O;
	wire [15:0] RMUX_T2_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T2_NORTH_B16_sel_inst0_O;
	wire [15:0] RMUX_T2_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T2_SOUTH_B16_sel_inst0_O;
	wire [15:0] RMUX_T2_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T2_WEST_B16_sel_inst0_O;
	wire [1:0] SB_T0_EAST_SB_OUT_B16_sel_inst0_O;
	wire [1:0] SB_T0_NORTH_SB_OUT_B16_sel_inst0_O;
	wire [1:0] SB_T0_SOUTH_SB_OUT_B16_sel_inst0_O;
	wire [1:0] SB_T0_WEST_SB_OUT_B16_sel_inst0_O;
	wire [1:0] SB_T1_EAST_SB_OUT_B16_sel_inst0_O;
	wire [1:0] SB_T1_NORTH_SB_OUT_B16_sel_inst0_O;
	wire [1:0] SB_T1_SOUTH_SB_OUT_B16_sel_inst0_O;
	wire [1:0] SB_T1_WEST_SB_OUT_B16_sel_inst0_O;
	wire [1:0] SB_T2_EAST_SB_OUT_B16_sel_inst0_O;
	wire [1:0] SB_T2_NORTH_SB_OUT_B16_sel_inst0_O;
	wire [1:0] SB_T2_SOUTH_SB_OUT_B16_sel_inst0_O;
	wire [1:0] SB_T2_WEST_SB_OUT_B16_sel_inst0_O;
	wire [15:0] WIRE_SB_T0_EAST_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T0_NORTH_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T0_SOUTH_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T0_WEST_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T1_EAST_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T1_NORTH_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T1_SOUTH_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T1_WEST_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T2_EAST_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T2_NORTH_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T2_SOUTH_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T2_WEST_SB_IN_B16_O;
	wire ZextWrapper_4_32_inst0$bit_const_0_None_out;
	wire [3:0] ZextWrapper_4_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_4_32_inst0$self_O_in;
	wire [0:0] and1_inst0_out;
	wire [0:0] and1_inst1_out;
	wire [0:0] and1_inst10_out;
	wire [0:0] and1_inst11_out;
	wire [0:0] and1_inst2_out;
	wire [0:0] and1_inst3_out;
	wire [0:0] and1_inst4_out;
	wire [0:0] and1_inst5_out;
	wire [0:0] and1_inst6_out;
	wire [0:0] and1_inst7_out;
	wire [0:0] and1_inst8_out;
	wire [0:0] and1_inst9_out;
	wire [31:0] config_reg_0_O;
	wire [3:0] config_reg_1_O;
	wire [0:0] const_1_1_out;
	wire coreir_eq_1_inst0_out;
	wire coreir_eq_1_inst1_out;
	wire coreir_eq_1_inst10_out;
	wire coreir_eq_1_inst11_out;
	wire coreir_eq_1_inst2_out;
	wire coreir_eq_1_inst3_out;
	wire coreir_eq_1_inst4_out;
	wire coreir_eq_1_inst5_out;
	wire coreir_eq_1_inst6_out;
	wire coreir_eq_1_inst7_out;
	wire coreir_eq_1_inst8_out;
	wire coreir_eq_1_inst9_out;
	coreir_not #(.width(1)) Invert1_inst0(
		.in(stall),
		.out(Invert1_inst0_out)
	);
	commonlib_muxn__N4__width16 MUX_SB_T0_EAST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0(
		.in_data_0(WIRE_SB_T0_WEST_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T2_NORTH_SB_IN_B16_O),
		.in_data_3(alu_res),
		.in_sel(SB_T0_EAST_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T0_EAST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out)
	);
	commonlib_muxn__N4__width16 MUX_SB_T0_NORTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0(
		.in_data_0(WIRE_SB_T0_WEST_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T1_EAST_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
		.in_data_3(alu_res),
		.in_sel(SB_T0_NORTH_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T0_NORTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out)
	);
	commonlib_muxn__N4__width16 MUX_SB_T0_SOUTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0(
		.in_data_0(WIRE_SB_T1_EAST_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T0_NORTH_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T1_WEST_SB_IN_B16_O),
		.in_data_3(alu_res),
		.in_sel(SB_T0_SOUTH_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T0_SOUTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out)
	);
	commonlib_muxn__N4__width16 MUX_SB_T0_WEST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0(
		.in_data_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
		.in_data_3(alu_res),
		.in_sel(SB_T0_WEST_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T0_WEST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out)
	);
	commonlib_muxn__N4__width16 MUX_SB_T1_EAST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0(
		.in_data_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T1_WEST_SB_IN_B16_O),
		.in_data_3(alu_res),
		.in_sel(SB_T1_EAST_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T1_EAST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out)
	);
	commonlib_muxn__N4__width16 MUX_SB_T1_NORTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0(
		.in_data_0(WIRE_SB_T2_EAST_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T2_WEST_SB_IN_B16_O),
		.in_data_3(alu_res),
		.in_sel(SB_T1_NORTH_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T1_NORTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out)
	);
	commonlib_muxn__N4__width16 MUX_SB_T1_SOUTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0(
		.in_data_0(WIRE_SB_T0_EAST_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T1_NORTH_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T2_WEST_SB_IN_B16_O),
		.in_data_3(alu_res),
		.in_sel(SB_T1_SOUTH_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T1_SOUTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out)
	);
	commonlib_muxn__N4__width16 MUX_SB_T1_WEST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0(
		.in_data_0(WIRE_SB_T2_NORTH_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T1_EAST_SB_IN_B16_O),
		.in_data_3(alu_res),
		.in_sel(SB_T1_WEST_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T1_WEST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out)
	);
	commonlib_muxn__N4__width16 MUX_SB_T2_EAST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0(
		.in_data_0(WIRE_SB_T1_NORTH_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T2_WEST_SB_IN_B16_O),
		.in_data_3(alu_res),
		.in_sel(SB_T2_EAST_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T2_EAST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out)
	);
	commonlib_muxn__N4__width16 MUX_SB_T2_NORTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0(
		.in_data_0(WIRE_SB_T1_WEST_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T0_EAST_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
		.in_data_3(alu_res),
		.in_sel(SB_T2_NORTH_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T2_NORTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out)
	);
	commonlib_muxn__N4__width16 MUX_SB_T2_SOUTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0(
		.in_data_0(WIRE_SB_T0_WEST_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T2_EAST_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T2_NORTH_SB_IN_B16_O),
		.in_data_3(alu_res),
		.in_sel(SB_T2_SOUTH_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T2_SOUTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out)
	);
	commonlib_muxn__N4__width16 MUX_SB_T2_WEST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0(
		.in_data_0(WIRE_SB_T1_NORTH_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T2_EAST_SB_IN_B16_O),
		.in_data_3(alu_res),
		.in_sel(SB_T2_WEST_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T2_WEST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out)
	);
	coreir_mux #(.width(32)) MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join(
		.in0(config_reg_0_O),
		.in1(ZextWrapper_4_32_inst0$self_O_in),
		.sel(config_config_addr[0]),
		.out(MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out)
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_EAST_B16(
		.I(MUX_SB_T0_EAST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.O(REG_T0_EAST_B16_O),
		.CLK(clk),
		.CE(and1_inst2_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_NORTH_B16(
		.I(MUX_SB_T0_NORTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.O(REG_T0_NORTH_B16_O),
		.CLK(clk),
		.CE(and1_inst0_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_SOUTH_B16(
		.I(MUX_SB_T0_SOUTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.O(REG_T0_SOUTH_B16_O),
		.CLK(clk),
		.CE(and1_inst1_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_WEST_B16(
		.I(MUX_SB_T0_WEST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.O(REG_T0_WEST_B16_O),
		.CLK(clk),
		.CE(and1_inst3_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_EAST_B16(
		.I(MUX_SB_T1_EAST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.O(REG_T1_EAST_B16_O),
		.CLK(clk),
		.CE(and1_inst6_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_NORTH_B16(
		.I(MUX_SB_T1_NORTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.O(REG_T1_NORTH_B16_O),
		.CLK(clk),
		.CE(and1_inst4_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_SOUTH_B16(
		.I(MUX_SB_T1_SOUTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.O(REG_T1_SOUTH_B16_O),
		.CLK(clk),
		.CE(and1_inst5_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_WEST_B16(
		.I(MUX_SB_T1_WEST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.O(REG_T1_WEST_B16_O),
		.CLK(clk),
		.CE(and1_inst7_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_EAST_B16(
		.I(MUX_SB_T2_EAST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.O(REG_T2_EAST_B16_O),
		.CLK(clk),
		.CE(and1_inst10_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_NORTH_B16(
		.I(MUX_SB_T2_NORTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.O(REG_T2_NORTH_B16_O),
		.CLK(clk),
		.CE(and1_inst8_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_SOUTH_B16(
		.I(MUX_SB_T2_SOUTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.O(REG_T2_SOUTH_B16_O),
		.CLK(clk),
		.CE(and1_inst9_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_WEST_B16(
		.I(MUX_SB_T2_WEST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.O(REG_T2_WEST_B16_O),
		.CLK(clk),
		.CE(and1_inst11_out[0])
	);
	coreir_mux #(.width(16)) RMUX_T0_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T0_EAST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.in1(REG_T0_EAST_B16_O),
		.sel(RMUX_T0_EAST_B16_sel_inst0_O[0]),
		.out(RMUX_T0_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T0_EAST_B16_sel RMUX_T0_EAST_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T0_EAST_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T0_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T0_NORTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.in1(REG_T0_NORTH_B16_O),
		.sel(RMUX_T0_NORTH_B16_sel_inst0_O[0]),
		.out(RMUX_T0_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T0_NORTH_B16_sel RMUX_T0_NORTH_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T0_NORTH_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T0_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T0_SOUTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.in1(REG_T0_SOUTH_B16_O),
		.sel(RMUX_T0_SOUTH_B16_sel_inst0_O[0]),
		.out(RMUX_T0_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T0_SOUTH_B16_sel RMUX_T0_SOUTH_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T0_SOUTH_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T0_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T0_WEST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.in1(REG_T0_WEST_B16_O),
		.sel(RMUX_T0_WEST_B16_sel_inst0_O[0]),
		.out(RMUX_T0_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T0_WEST_B16_sel RMUX_T0_WEST_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T0_WEST_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T1_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T1_EAST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.in1(REG_T1_EAST_B16_O),
		.sel(RMUX_T1_EAST_B16_sel_inst0_O[0]),
		.out(RMUX_T1_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T1_EAST_B16_sel RMUX_T1_EAST_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T1_EAST_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T1_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T1_NORTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.in1(REG_T1_NORTH_B16_O),
		.sel(RMUX_T1_NORTH_B16_sel_inst0_O[0]),
		.out(RMUX_T1_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T1_NORTH_B16_sel RMUX_T1_NORTH_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T1_NORTH_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T1_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T1_SOUTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.in1(REG_T1_SOUTH_B16_O),
		.sel(RMUX_T1_SOUTH_B16_sel_inst0_O[0]),
		.out(RMUX_T1_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T1_SOUTH_B16_sel RMUX_T1_SOUTH_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T1_SOUTH_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T1_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T1_WEST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.in1(REG_T1_WEST_B16_O),
		.sel(RMUX_T1_WEST_B16_sel_inst0_O[0]),
		.out(RMUX_T1_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T1_WEST_B16_sel RMUX_T1_WEST_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T1_WEST_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T2_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T2_EAST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.in1(REG_T2_EAST_B16_O),
		.sel(RMUX_T2_EAST_B16_sel_inst0_O[0]),
		.out(RMUX_T2_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T2_EAST_B16_sel RMUX_T2_EAST_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T2_EAST_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T2_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T2_NORTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.in1(REG_T2_NORTH_B16_O),
		.sel(RMUX_T2_NORTH_B16_sel_inst0_O[0]),
		.out(RMUX_T2_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T2_NORTH_B16_sel RMUX_T2_NORTH_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T2_NORTH_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T2_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T2_SOUTH_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.in1(REG_T2_SOUTH_B16_O),
		.sel(RMUX_T2_SOUTH_B16_sel_inst0_O[0]),
		.out(RMUX_T2_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T2_SOUTH_B16_sel RMUX_T2_SOUTH_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T2_SOUTH_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T2_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T2_WEST_SB_OUT_B16$Mux4xBits16_inst0$coreir_commonlib_mux4x16_inst0_out),
		.in1(REG_T2_WEST_B16_O),
		.sel(RMUX_T2_WEST_B16_sel_inst0_O[0]),
		.out(RMUX_T2_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T2_WEST_B16_sel RMUX_T2_WEST_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T2_WEST_B16_sel_inst0_O)
	);
	SB_T0_EAST_SB_OUT_B16_sel SB_T0_EAST_SB_OUT_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T0_EAST_SB_OUT_B16_sel_inst0_O)
	);
	SB_T0_NORTH_SB_OUT_B16_sel SB_T0_NORTH_SB_OUT_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T0_NORTH_SB_OUT_B16_sel_inst0_O)
	);
	SB_T0_SOUTH_SB_OUT_B16_sel SB_T0_SOUTH_SB_OUT_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T0_SOUTH_SB_OUT_B16_sel_inst0_O)
	);
	SB_T0_WEST_SB_OUT_B16_sel SB_T0_WEST_SB_OUT_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T0_WEST_SB_OUT_B16_sel_inst0_O)
	);
	SB_T1_EAST_SB_OUT_B16_sel SB_T1_EAST_SB_OUT_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T1_EAST_SB_OUT_B16_sel_inst0_O)
	);
	SB_T1_NORTH_SB_OUT_B16_sel SB_T1_NORTH_SB_OUT_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T1_NORTH_SB_OUT_B16_sel_inst0_O)
	);
	SB_T1_SOUTH_SB_OUT_B16_sel SB_T1_SOUTH_SB_OUT_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T1_SOUTH_SB_OUT_B16_sel_inst0_O)
	);
	SB_T1_WEST_SB_OUT_B16_sel SB_T1_WEST_SB_OUT_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T1_WEST_SB_OUT_B16_sel_inst0_O)
	);
	SB_T2_EAST_SB_OUT_B16_sel SB_T2_EAST_SB_OUT_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T2_EAST_SB_OUT_B16_sel_inst0_O)
	);
	SB_T2_NORTH_SB_OUT_B16_sel SB_T2_NORTH_SB_OUT_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T2_NORTH_SB_OUT_B16_sel_inst0_O)
	);
	SB_T2_SOUTH_SB_OUT_B16_sel SB_T2_SOUTH_SB_OUT_B16_sel_inst0(
		.I(config_reg_1_O),
		.O(SB_T2_SOUTH_SB_OUT_B16_sel_inst0_O)
	);
	SB_T2_WEST_SB_OUT_B16_sel SB_T2_WEST_SB_OUT_B16_sel_inst0(
		.I(config_reg_1_O),
		.O(SB_T2_WEST_SB_OUT_B16_sel_inst0_O)
	);
	MuxWrapper_1_16 WIRE_SB_T0_EAST_SB_IN_B16(
		.I(SB_T0_EAST_SB_IN_B16),
		.O(WIRE_SB_T0_EAST_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T0_NORTH_SB_IN_B16(
		.I(SB_T0_NORTH_SB_IN_B16),
		.O(WIRE_SB_T0_NORTH_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T0_SOUTH_SB_IN_B16(
		.I(SB_T0_SOUTH_SB_IN_B16),
		.O(WIRE_SB_T0_SOUTH_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T0_WEST_SB_IN_B16(
		.I(SB_T0_WEST_SB_IN_B16),
		.O(WIRE_SB_T0_WEST_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T1_EAST_SB_IN_B16(
		.I(SB_T1_EAST_SB_IN_B16),
		.O(WIRE_SB_T1_EAST_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T1_NORTH_SB_IN_B16(
		.I(SB_T1_NORTH_SB_IN_B16),
		.O(WIRE_SB_T1_NORTH_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T1_SOUTH_SB_IN_B16(
		.I(SB_T1_SOUTH_SB_IN_B16),
		.O(WIRE_SB_T1_SOUTH_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T1_WEST_SB_IN_B16(
		.I(SB_T1_WEST_SB_IN_B16),
		.O(WIRE_SB_T1_WEST_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T2_EAST_SB_IN_B16(
		.I(SB_T2_EAST_SB_IN_B16),
		.O(WIRE_SB_T2_EAST_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T2_NORTH_SB_IN_B16(
		.I(SB_T2_NORTH_SB_IN_B16),
		.O(WIRE_SB_T2_NORTH_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T2_SOUTH_SB_IN_B16(
		.I(SB_T2_SOUTH_SB_IN_B16),
		.O(WIRE_SB_T2_SOUTH_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T2_WEST_SB_IN_B16(
		.I(SB_T2_WEST_SB_IN_B16),
		.O(WIRE_SB_T2_WEST_SB_IN_B16_O)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_4_32_inst0$bit_const_0_None(.out(ZextWrapper_4_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit4 ZextWrapper_4_32_inst0$self_I(
		.in(config_reg_1_O),
		.out(ZextWrapper_4_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_4_32_inst0$self_O_out;
	assign ZextWrapper_4_32_inst0$self_O_out = {ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$self_I_out[3:0]};
	mantle_wire__typeBitIn32 ZextWrapper_4_32_inst0$self_O(
		.in(ZextWrapper_4_32_inst0$self_O_in),
		.out(ZextWrapper_4_32_inst0$self_O_out)
	);
	coreir_and #(.width(1)) and1_inst0(
		.in0(coreir_eq_1_inst0_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst0_out)
	);
	coreir_and #(.width(1)) and1_inst1(
		.in0(coreir_eq_1_inst1_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst1_out)
	);
	coreir_and #(.width(1)) and1_inst10(
		.in0(coreir_eq_1_inst10_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst10_out)
	);
	coreir_and #(.width(1)) and1_inst11(
		.in0(coreir_eq_1_inst11_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst11_out)
	);
	coreir_and #(.width(1)) and1_inst2(
		.in0(coreir_eq_1_inst2_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst2_out)
	);
	coreir_and #(.width(1)) and1_inst3(
		.in0(coreir_eq_1_inst3_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst3_out)
	);
	coreir_and #(.width(1)) and1_inst4(
		.in0(coreir_eq_1_inst4_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst4_out)
	);
	coreir_and #(.width(1)) and1_inst5(
		.in0(coreir_eq_1_inst5_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst5_out)
	);
	coreir_and #(.width(1)) and1_inst6(
		.in0(coreir_eq_1_inst6_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst6_out)
	);
	coreir_and #(.width(1)) and1_inst7(
		.in0(coreir_eq_1_inst7_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst7_out)
	);
	coreir_and #(.width(1)) and1_inst8(
		.in0(coreir_eq_1_inst8_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst8_out)
	);
	coreir_and #(.width(1)) and1_inst9(
		.in0(coreir_eq_1_inst9_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst9_out)
	);
	ConfigRegister_32_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_4_8_32_1 config_reg_1(
		.clk(clk),
		.reset(reset),
		.O(config_reg_1_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	coreir_const #(
		.value(1'h1),
		.width(1)
	) const_1_1(.out(const_1_1_out));
	coreir_eq #(.width(1)) coreir_eq_1_inst0(
		.in0(const_1_1_out),
		.in1(RMUX_T0_NORTH_B16_sel_inst0_O),
		.out(coreir_eq_1_inst0_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst1(
		.in0(const_1_1_out),
		.in1(RMUX_T0_SOUTH_B16_sel_inst0_O),
		.out(coreir_eq_1_inst1_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst10(
		.in0(const_1_1_out),
		.in1(RMUX_T2_EAST_B16_sel_inst0_O),
		.out(coreir_eq_1_inst10_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst11(
		.in0(const_1_1_out),
		.in1(RMUX_T2_WEST_B16_sel_inst0_O),
		.out(coreir_eq_1_inst11_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst2(
		.in0(const_1_1_out),
		.in1(RMUX_T0_EAST_B16_sel_inst0_O),
		.out(coreir_eq_1_inst2_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst3(
		.in0(const_1_1_out),
		.in1(RMUX_T0_WEST_B16_sel_inst0_O),
		.out(coreir_eq_1_inst3_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst4(
		.in0(const_1_1_out),
		.in1(RMUX_T1_NORTH_B16_sel_inst0_O),
		.out(coreir_eq_1_inst4_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst5(
		.in0(const_1_1_out),
		.in1(RMUX_T1_SOUTH_B16_sel_inst0_O),
		.out(coreir_eq_1_inst5_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst6(
		.in0(const_1_1_out),
		.in1(RMUX_T1_EAST_B16_sel_inst0_O),
		.out(coreir_eq_1_inst6_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst7(
		.in0(const_1_1_out),
		.in1(RMUX_T1_WEST_B16_sel_inst0_O),
		.out(coreir_eq_1_inst7_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst8(
		.in0(const_1_1_out),
		.in1(RMUX_T2_NORTH_B16_sel_inst0_O),
		.out(coreir_eq_1_inst8_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst9(
		.in0(const_1_1_out),
		.in1(RMUX_T2_SOUTH_B16_sel_inst0_O),
		.out(coreir_eq_1_inst9_out)
	);
	assign SB_T0_EAST_SB_OUT_B16 = RMUX_T0_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T0_NORTH_SB_OUT_B16 = RMUX_T0_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T0_SOUTH_SB_OUT_B16 = RMUX_T0_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T0_WEST_SB_OUT_B16 = RMUX_T0_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T1_EAST_SB_OUT_B16 = RMUX_T1_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T1_NORTH_SB_OUT_B16 = RMUX_T1_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T1_SOUTH_SB_OUT_B16 = RMUX_T1_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T1_WEST_SB_OUT_B16 = RMUX_T1_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T2_EAST_SB_OUT_B16 = RMUX_T2_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T2_NORTH_SB_OUT_B16 = RMUX_T2_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T2_SOUTH_SB_OUT_B16 = RMUX_T2_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T2_WEST_SB_OUT_B16 = RMUX_T2_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign read_config_data = MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
endmodule
module ConfigRegister_30_8_32_0 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [29:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [29:0] Register_inst0_O;
	wire [7:0] const_0_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq10 Register_inst0(
		.I(config_data[29:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h00),
		.width(8)
	) const_0_8(.out(const_0_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_0_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_28_8_32_48 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [27:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [27:0] Register_inst0_O;
	wire [7:0] const_48_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq8 Register_inst0(
		.I(config_data[27:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h30),
		.width(8)
	) const_48_8(.out(const_48_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_48_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_26_8_32_0 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [25:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [25:0] Register_inst0_O;
	wire [7:0] const_0_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq4 Register_inst0(
		.I(config_data[25:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h00),
		.width(8)
	) const_0_8(.out(const_0_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_0_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_25_8_32_71 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [24:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [24:0] Register_inst0_O;
	wire [7:0] const_71_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq7 Register_inst0(
		.I(config_data[24:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h47),
		.width(8)
	) const_71_8(.out(const_71_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_71_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_25_8_32_41 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [24:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [24:0] Register_inst0_O;
	wire [7:0] const_41_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq7 Register_inst0(
		.I(config_data[24:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h29),
		.width(8)
	) const_41_8(.out(const_41_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_41_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_20_8_32_66 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [19:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [19:0] Register_inst0_O;
	wire [7:0] const_66_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq6 Register_inst0(
		.I(config_data[19:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h42),
		.width(8)
	) const_66_8(.out(const_66_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_66_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_20_8_32_63 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [19:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [19:0] Register_inst0_O;
	wire [7:0] const_63_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq6 Register_inst0(
		.I(config_data[19:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h3f),
		.width(8)
	) const_63_8(.out(const_63_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_63_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_20_8_32_51 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [19:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [19:0] Register_inst0_O;
	wire [7:0] const_51_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq6 Register_inst0(
		.I(config_data[19:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h33),
		.width(8)
	) const_51_8(.out(const_51_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_51_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_20_8_32_37 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [19:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [19:0] Register_inst0_O;
	wire [7:0] const_37_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq6 Register_inst0(
		.I(config_data[19:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h25),
		.width(8)
	) const_37_8(.out(const_37_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_37_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_20_8_32_34 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [19:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [19:0] Register_inst0_O;
	wire [7:0] const_34_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq6 Register_inst0(
		.I(config_data[19:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h22),
		.width(8)
	) const_34_8(.out(const_34_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_34_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_20_8_32_22 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [19:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [19:0] Register_inst0_O;
	wire [7:0] const_22_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq6 Register_inst0(
		.I(config_data[19:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h16),
		.width(8)
	) const_22_8(.out(const_22_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_22_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_20_8_32_19 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [19:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [19:0] Register_inst0_O;
	wire [7:0] const_19_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq6 Register_inst0(
		.I(config_data[19:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h13),
		.width(8)
	) const_19_8(.out(const_19_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_19_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_18_8_32_1 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [17:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [17:0] Register_inst0_O;
	wire [7:0] const_1_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq11 Register_inst0(
		.I(config_data[17:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h01),
		.width(8)
	) const_1_8(.out(const_1_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_1_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module SB_ID0_3TRACKS_B1_MemCore (
	SB_T0_EAST_SB_IN_B1,
	SB_T0_EAST_SB_OUT_B1,
	SB_T0_NORTH_SB_IN_B1,
	SB_T0_NORTH_SB_OUT_B1,
	SB_T0_SOUTH_SB_IN_B1,
	SB_T0_SOUTH_SB_OUT_B1,
	SB_T0_WEST_SB_IN_B1,
	SB_T0_WEST_SB_OUT_B1,
	SB_T1_EAST_SB_IN_B1,
	SB_T1_EAST_SB_OUT_B1,
	SB_T1_NORTH_SB_IN_B1,
	SB_T1_NORTH_SB_OUT_B1,
	SB_T1_SOUTH_SB_IN_B1,
	SB_T1_SOUTH_SB_OUT_B1,
	SB_T1_WEST_SB_IN_B1,
	SB_T1_WEST_SB_OUT_B1,
	SB_T2_EAST_SB_IN_B1,
	SB_T2_EAST_SB_OUT_B1,
	SB_T2_NORTH_SB_IN_B1,
	SB_T2_NORTH_SB_OUT_B1,
	SB_T2_SOUTH_SB_IN_B1,
	SB_T2_SOUTH_SB_OUT_B1,
	SB_T2_WEST_SB_IN_B1,
	SB_T2_WEST_SB_OUT_B1,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	output_width_1_num_0,
	output_width_1_num_1,
	output_width_1_num_2,
	read_config_data,
	reset,
	stall
);
	input [0:0] SB_T0_EAST_SB_IN_B1;
	output [0:0] SB_T0_EAST_SB_OUT_B1;
	input [0:0] SB_T0_NORTH_SB_IN_B1;
	output [0:0] SB_T0_NORTH_SB_OUT_B1;
	input [0:0] SB_T0_SOUTH_SB_IN_B1;
	output [0:0] SB_T0_SOUTH_SB_OUT_B1;
	input [0:0] SB_T0_WEST_SB_IN_B1;
	output [0:0] SB_T0_WEST_SB_OUT_B1;
	input [0:0] SB_T1_EAST_SB_IN_B1;
	output [0:0] SB_T1_EAST_SB_OUT_B1;
	input [0:0] SB_T1_NORTH_SB_IN_B1;
	output [0:0] SB_T1_NORTH_SB_OUT_B1;
	input [0:0] SB_T1_SOUTH_SB_IN_B1;
	output [0:0] SB_T1_SOUTH_SB_OUT_B1;
	input [0:0] SB_T1_WEST_SB_IN_B1;
	output [0:0] SB_T1_WEST_SB_OUT_B1;
	input [0:0] SB_T2_EAST_SB_IN_B1;
	output [0:0] SB_T2_EAST_SB_OUT_B1;
	input [0:0] SB_T2_NORTH_SB_IN_B1;
	output [0:0] SB_T2_NORTH_SB_OUT_B1;
	input [0:0] SB_T2_SOUTH_SB_IN_B1;
	output [0:0] SB_T2_SOUTH_SB_OUT_B1;
	input [0:0] SB_T2_WEST_SB_IN_B1;
	output [0:0] SB_T2_WEST_SB_OUT_B1;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	input [0:0] output_width_1_num_0;
	input [0:0] output_width_1_num_1;
	input [0:0] output_width_1_num_2;
	output [31:0] read_config_data;
	input reset;
	input [0:0] stall;
	wire [0:0] Invert1_inst0_out;
	wire [0:0] MUX_SB_T0_EAST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out;
	wire [0:0] MUX_SB_T0_NORTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out;
	wire [0:0] MUX_SB_T0_SOUTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out;
	wire [0:0] MUX_SB_T0_WEST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out;
	wire [0:0] MUX_SB_T1_EAST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out;
	wire [0:0] MUX_SB_T1_NORTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out;
	wire [0:0] MUX_SB_T1_SOUTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out;
	wire [0:0] MUX_SB_T1_WEST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out;
	wire [0:0] MUX_SB_T2_EAST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out;
	wire [0:0] MUX_SB_T2_NORTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out;
	wire [0:0] MUX_SB_T2_SOUTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out;
	wire [0:0] MUX_SB_T2_WEST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out;
	wire [31:0] MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
	wire [0:0] REG_T0_EAST_B1_O;
	wire [0:0] REG_T0_NORTH_B1_O;
	wire [0:0] REG_T0_SOUTH_B1_O;
	wire [0:0] REG_T0_WEST_B1_O;
	wire [0:0] REG_T1_EAST_B1_O;
	wire [0:0] REG_T1_NORTH_B1_O;
	wire [0:0] REG_T1_SOUTH_B1_O;
	wire [0:0] REG_T1_WEST_B1_O;
	wire [0:0] REG_T2_EAST_B1_O;
	wire [0:0] REG_T2_NORTH_B1_O;
	wire [0:0] REG_T2_SOUTH_B1_O;
	wire [0:0] REG_T2_WEST_B1_O;
	wire [0:0] RMUX_T0_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T0_EAST_B1_sel_inst0_O;
	wire [0:0] RMUX_T0_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T0_NORTH_B1_sel_inst0_O;
	wire [0:0] RMUX_T0_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T0_SOUTH_B1_sel_inst0_O;
	wire [0:0] RMUX_T0_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T0_WEST_B1_sel_inst0_O;
	wire [0:0] RMUX_T1_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T1_EAST_B1_sel_inst0_O;
	wire [0:0] RMUX_T1_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T1_NORTH_B1_sel_inst0_O;
	wire [0:0] RMUX_T1_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T1_SOUTH_B1_sel_inst0_O;
	wire [0:0] RMUX_T1_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T1_WEST_B1_sel_inst0_O;
	wire [0:0] RMUX_T2_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T2_EAST_B1_sel_inst0_O;
	wire [0:0] RMUX_T2_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T2_NORTH_B1_sel_inst0_O;
	wire [0:0] RMUX_T2_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T2_SOUTH_B1_sel_inst0_O;
	wire [0:0] RMUX_T2_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] RMUX_T2_WEST_B1_sel_inst0_O;
	wire [2:0] SB_T0_EAST_SB_OUT_B1_sel_inst0_O;
	wire [2:0] SB_T0_NORTH_SB_OUT_B1_sel_inst0_O;
	wire [2:0] SB_T0_SOUTH_SB_OUT_B1_sel_inst0_O;
	wire [2:0] SB_T0_WEST_SB_OUT_B1_sel_inst0_O;
	wire [2:0] SB_T1_EAST_SB_OUT_B1_sel_inst0_O;
	wire [2:0] SB_T1_NORTH_SB_OUT_B1_sel_inst0_O;
	wire [2:0] SB_T1_SOUTH_SB_OUT_B1_sel_inst0_O;
	wire [2:0] SB_T1_WEST_SB_OUT_B1_sel_inst0_O;
	wire [2:0] SB_T2_EAST_SB_OUT_B1_sel_inst0_O;
	wire [2:0] SB_T2_NORTH_SB_OUT_B1_sel_inst0_O;
	wire [2:0] SB_T2_SOUTH_SB_OUT_B1_sel_inst0_O;
	wire [2:0] SB_T2_WEST_SB_OUT_B1_sel_inst0_O;
	wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1_O;
	wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1_O;
	wire ZextWrapper_18_32_inst0$bit_const_0_None_out;
	wire [17:0] ZextWrapper_18_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_18_32_inst0$self_O_in;
	wire ZextWrapper_30_32_inst0$bit_const_0_None_out;
	wire [29:0] ZextWrapper_30_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_30_32_inst0$self_O_in;
	wire [0:0] and1_inst0_out;
	wire [0:0] and1_inst1_out;
	wire [0:0] and1_inst10_out;
	wire [0:0] and1_inst11_out;
	wire [0:0] and1_inst2_out;
	wire [0:0] and1_inst3_out;
	wire [0:0] and1_inst4_out;
	wire [0:0] and1_inst5_out;
	wire [0:0] and1_inst6_out;
	wire [0:0] and1_inst7_out;
	wire [0:0] and1_inst8_out;
	wire [0:0] and1_inst9_out;
	wire [29:0] config_reg_0_O;
	wire [17:0] config_reg_1_O;
	wire [0:0] const_1_1_out;
	wire coreir_eq_1_inst0_out;
	wire coreir_eq_1_inst1_out;
	wire coreir_eq_1_inst10_out;
	wire coreir_eq_1_inst11_out;
	wire coreir_eq_1_inst2_out;
	wire coreir_eq_1_inst3_out;
	wire coreir_eq_1_inst4_out;
	wire coreir_eq_1_inst5_out;
	wire coreir_eq_1_inst6_out;
	wire coreir_eq_1_inst7_out;
	wire coreir_eq_1_inst8_out;
	wire coreir_eq_1_inst9_out;
	coreir_not #(.width(1)) Invert1_inst0(
		.in(stall),
		.out(Invert1_inst0_out)
	);
	commonlib_muxn__N6__width1 MUX_SB_T0_EAST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0(
		.in_data_0(WIRE_SB_T0_WEST_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T2_NORTH_SB_IN_B1_O),
		.in_data_3(output_width_1_num_0),
		.in_data_4(output_width_1_num_1),
		.in_data_5(output_width_1_num_2),
		.in_sel(SB_T0_EAST_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T0_EAST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out)
	);
	commonlib_muxn__N6__width1 MUX_SB_T0_NORTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0(
		.in_data_0(WIRE_SB_T0_WEST_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T1_EAST_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
		.in_data_3(output_width_1_num_0),
		.in_data_4(output_width_1_num_1),
		.in_data_5(output_width_1_num_2),
		.in_sel(SB_T0_NORTH_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T0_NORTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out)
	);
	commonlib_muxn__N6__width1 MUX_SB_T0_SOUTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0(
		.in_data_0(WIRE_SB_T1_EAST_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T0_NORTH_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T1_WEST_SB_IN_B1_O),
		.in_data_3(output_width_1_num_0),
		.in_data_4(output_width_1_num_1),
		.in_data_5(output_width_1_num_2),
		.in_sel(SB_T0_SOUTH_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T0_SOUTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out)
	);
	commonlib_muxn__N6__width1 MUX_SB_T0_WEST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0(
		.in_data_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
		.in_data_3(output_width_1_num_0),
		.in_data_4(output_width_1_num_1),
		.in_data_5(output_width_1_num_2),
		.in_sel(SB_T0_WEST_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T0_WEST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out)
	);
	commonlib_muxn__N6__width1 MUX_SB_T1_EAST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0(
		.in_data_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T1_WEST_SB_IN_B1_O),
		.in_data_3(output_width_1_num_0),
		.in_data_4(output_width_1_num_1),
		.in_data_5(output_width_1_num_2),
		.in_sel(SB_T1_EAST_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T1_EAST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out)
	);
	commonlib_muxn__N6__width1 MUX_SB_T1_NORTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0(
		.in_data_0(WIRE_SB_T2_EAST_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T2_WEST_SB_IN_B1_O),
		.in_data_3(output_width_1_num_0),
		.in_data_4(output_width_1_num_1),
		.in_data_5(output_width_1_num_2),
		.in_sel(SB_T1_NORTH_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T1_NORTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out)
	);
	commonlib_muxn__N6__width1 MUX_SB_T1_SOUTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0(
		.in_data_0(WIRE_SB_T0_EAST_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T1_NORTH_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T2_WEST_SB_IN_B1_O),
		.in_data_3(output_width_1_num_0),
		.in_data_4(output_width_1_num_1),
		.in_data_5(output_width_1_num_2),
		.in_sel(SB_T1_SOUTH_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T1_SOUTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out)
	);
	commonlib_muxn__N6__width1 MUX_SB_T1_WEST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0(
		.in_data_0(WIRE_SB_T2_NORTH_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T1_EAST_SB_IN_B1_O),
		.in_data_3(output_width_1_num_0),
		.in_data_4(output_width_1_num_1),
		.in_data_5(output_width_1_num_2),
		.in_sel(SB_T1_WEST_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T1_WEST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out)
	);
	commonlib_muxn__N6__width1 MUX_SB_T2_EAST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0(
		.in_data_0(WIRE_SB_T1_NORTH_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T2_WEST_SB_IN_B1_O),
		.in_data_3(output_width_1_num_0),
		.in_data_4(output_width_1_num_1),
		.in_data_5(output_width_1_num_2),
		.in_sel(SB_T2_EAST_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T2_EAST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out)
	);
	commonlib_muxn__N6__width1 MUX_SB_T2_NORTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0(
		.in_data_0(WIRE_SB_T1_WEST_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T0_EAST_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
		.in_data_3(output_width_1_num_0),
		.in_data_4(output_width_1_num_1),
		.in_data_5(output_width_1_num_2),
		.in_sel(SB_T2_NORTH_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T2_NORTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out)
	);
	commonlib_muxn__N6__width1 MUX_SB_T2_SOUTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0(
		.in_data_0(WIRE_SB_T0_WEST_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T2_EAST_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T2_NORTH_SB_IN_B1_O),
		.in_data_3(output_width_1_num_0),
		.in_data_4(output_width_1_num_1),
		.in_data_5(output_width_1_num_2),
		.in_sel(SB_T2_SOUTH_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T2_SOUTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out)
	);
	commonlib_muxn__N6__width1 MUX_SB_T2_WEST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0(
		.in_data_0(WIRE_SB_T1_NORTH_SB_IN_B1_O),
		.in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
		.in_data_2(WIRE_SB_T2_EAST_SB_IN_B1_O),
		.in_data_3(output_width_1_num_0),
		.in_data_4(output_width_1_num_1),
		.in_data_5(output_width_1_num_2),
		.in_sel(SB_T2_WEST_SB_OUT_B1_sel_inst0_O),
		.out(MUX_SB_T2_WEST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out)
	);
	coreir_mux #(.width(32)) MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join(
		.in0(ZextWrapper_30_32_inst0$self_O_in),
		.in1(ZextWrapper_18_32_inst0$self_O_in),
		.sel(config_config_addr[0]),
		.out(MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out)
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_EAST_B1(
		.I(MUX_SB_T0_EAST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.O(REG_T0_EAST_B1_O),
		.CLK(clk),
		.CE(and1_inst2_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_NORTH_B1(
		.I(MUX_SB_T0_NORTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.O(REG_T0_NORTH_B1_O),
		.CLK(clk),
		.CE(and1_inst0_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_SOUTH_B1(
		.I(MUX_SB_T0_SOUTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.O(REG_T0_SOUTH_B1_O),
		.CLK(clk),
		.CE(and1_inst1_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_WEST_B1(
		.I(MUX_SB_T0_WEST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.O(REG_T0_WEST_B1_O),
		.CLK(clk),
		.CE(and1_inst3_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_EAST_B1(
		.I(MUX_SB_T1_EAST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.O(REG_T1_EAST_B1_O),
		.CLK(clk),
		.CE(and1_inst6_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_NORTH_B1(
		.I(MUX_SB_T1_NORTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.O(REG_T1_NORTH_B1_O),
		.CLK(clk),
		.CE(and1_inst4_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_SOUTH_B1(
		.I(MUX_SB_T1_SOUTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.O(REG_T1_SOUTH_B1_O),
		.CLK(clk),
		.CE(and1_inst5_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_WEST_B1(
		.I(MUX_SB_T1_WEST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.O(REG_T1_WEST_B1_O),
		.CLK(clk),
		.CE(and1_inst7_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_EAST_B1(
		.I(MUX_SB_T2_EAST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.O(REG_T2_EAST_B1_O),
		.CLK(clk),
		.CE(and1_inst10_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_NORTH_B1(
		.I(MUX_SB_T2_NORTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.O(REG_T2_NORTH_B1_O),
		.CLK(clk),
		.CE(and1_inst8_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_SOUTH_B1(
		.I(MUX_SB_T2_SOUTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.O(REG_T2_SOUTH_B1_O),
		.CLK(clk),
		.CE(and1_inst9_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_WEST_B1(
		.I(MUX_SB_T2_WEST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.O(REG_T2_WEST_B1_O),
		.CLK(clk),
		.CE(and1_inst11_out[0])
	);
	coreir_mux #(.width(1)) RMUX_T0_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T0_EAST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.in1(REG_T0_EAST_B1_O),
		.sel(RMUX_T0_EAST_B1_sel_inst0_O[0]),
		.out(RMUX_T0_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T0_EAST_B1_sel_unq1 RMUX_T0_EAST_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T0_EAST_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T0_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T0_NORTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.in1(REG_T0_NORTH_B1_O),
		.sel(RMUX_T0_NORTH_B1_sel_inst0_O[0]),
		.out(RMUX_T0_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T0_NORTH_B1_sel_unq1 RMUX_T0_NORTH_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T0_NORTH_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T0_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T0_SOUTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.in1(REG_T0_SOUTH_B1_O),
		.sel(RMUX_T0_SOUTH_B1_sel_inst0_O[0]),
		.out(RMUX_T0_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T0_SOUTH_B1_sel_unq1 RMUX_T0_SOUTH_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T0_SOUTH_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T0_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T0_WEST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.in1(REG_T0_WEST_B1_O),
		.sel(RMUX_T0_WEST_B1_sel_inst0_O[0]),
		.out(RMUX_T0_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T0_WEST_B1_sel_unq1 RMUX_T0_WEST_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T0_WEST_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T1_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T1_EAST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.in1(REG_T1_EAST_B1_O),
		.sel(RMUX_T1_EAST_B1_sel_inst0_O[0]),
		.out(RMUX_T1_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T1_EAST_B1_sel_unq1 RMUX_T1_EAST_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T1_EAST_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T1_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T1_NORTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.in1(REG_T1_NORTH_B1_O),
		.sel(RMUX_T1_NORTH_B1_sel_inst0_O[0]),
		.out(RMUX_T1_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T1_NORTH_B1_sel_unq1 RMUX_T1_NORTH_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T1_NORTH_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T1_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T1_SOUTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.in1(REG_T1_SOUTH_B1_O),
		.sel(RMUX_T1_SOUTH_B1_sel_inst0_O[0]),
		.out(RMUX_T1_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T1_SOUTH_B1_sel_unq1 RMUX_T1_SOUTH_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T1_SOUTH_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T1_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T1_WEST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.in1(REG_T1_WEST_B1_O),
		.sel(RMUX_T1_WEST_B1_sel_inst0_O[0]),
		.out(RMUX_T1_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T1_WEST_B1_sel_unq1 RMUX_T1_WEST_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T1_WEST_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T2_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T2_EAST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.in1(REG_T2_EAST_B1_O),
		.sel(RMUX_T2_EAST_B1_sel_inst0_O[0]),
		.out(RMUX_T2_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T2_EAST_B1_sel_unq1 RMUX_T2_EAST_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T2_EAST_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T2_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T2_NORTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.in1(REG_T2_NORTH_B1_O),
		.sel(RMUX_T2_NORTH_B1_sel_inst0_O[0]),
		.out(RMUX_T2_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T2_NORTH_B1_sel_unq1 RMUX_T2_NORTH_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T2_NORTH_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T2_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T2_SOUTH_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.in1(REG_T2_SOUTH_B1_O),
		.sel(RMUX_T2_SOUTH_B1_sel_inst0_O[0]),
		.out(RMUX_T2_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T2_SOUTH_B1_sel_unq1 RMUX_T2_SOUTH_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T2_SOUTH_B1_sel_inst0_O)
	);
	coreir_mux #(.width(1)) RMUX_T2_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(MUX_SB_T2_WEST_SB_OUT_B1$Mux6xBits1_inst0$coreir_commonlib_mux6x1_inst0_out),
		.in1(REG_T2_WEST_B1_O),
		.sel(RMUX_T2_WEST_B1_sel_inst0_O[0]),
		.out(RMUX_T2_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	RMUX_T2_WEST_B1_sel_unq1 RMUX_T2_WEST_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T2_WEST_B1_sel_inst0_O)
	);
	SB_T0_EAST_SB_OUT_B1_sel_unq1 SB_T0_EAST_SB_OUT_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T0_EAST_SB_OUT_B1_sel_inst0_O)
	);
	SB_T0_NORTH_SB_OUT_B1_sel_unq1 SB_T0_NORTH_SB_OUT_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T0_NORTH_SB_OUT_B1_sel_inst0_O)
	);
	SB_T0_SOUTH_SB_OUT_B1_sel_unq1 SB_T0_SOUTH_SB_OUT_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T0_SOUTH_SB_OUT_B1_sel_inst0_O)
	);
	SB_T0_WEST_SB_OUT_B1_sel_unq1 SB_T0_WEST_SB_OUT_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T0_WEST_SB_OUT_B1_sel_inst0_O)
	);
	SB_T1_EAST_SB_OUT_B1_sel_unq1 SB_T1_EAST_SB_OUT_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T1_EAST_SB_OUT_B1_sel_inst0_O)
	);
	SB_T1_NORTH_SB_OUT_B1_sel_unq1 SB_T1_NORTH_SB_OUT_B1_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T1_NORTH_SB_OUT_B1_sel_inst0_O)
	);
	SB_T1_SOUTH_SB_OUT_B1_sel_unq1 SB_T1_SOUTH_SB_OUT_B1_sel_inst0(
		.I(config_reg_1_O),
		.O(SB_T1_SOUTH_SB_OUT_B1_sel_inst0_O)
	);
	SB_T1_WEST_SB_OUT_B1_sel_unq1 SB_T1_WEST_SB_OUT_B1_sel_inst0(
		.I(config_reg_1_O),
		.O(SB_T1_WEST_SB_OUT_B1_sel_inst0_O)
	);
	SB_T2_EAST_SB_OUT_B1_sel_unq1 SB_T2_EAST_SB_OUT_B1_sel_inst0(
		.I(config_reg_1_O),
		.O(SB_T2_EAST_SB_OUT_B1_sel_inst0_O)
	);
	SB_T2_NORTH_SB_OUT_B1_sel_unq1 SB_T2_NORTH_SB_OUT_B1_sel_inst0(
		.I(config_reg_1_O),
		.O(SB_T2_NORTH_SB_OUT_B1_sel_inst0_O)
	);
	SB_T2_SOUTH_SB_OUT_B1_sel_unq1 SB_T2_SOUTH_SB_OUT_B1_sel_inst0(
		.I(config_reg_1_O),
		.O(SB_T2_SOUTH_SB_OUT_B1_sel_inst0_O)
	);
	SB_T2_WEST_SB_OUT_B1_sel_unq1 SB_T2_WEST_SB_OUT_B1_sel_inst0(
		.I(config_reg_1_O),
		.O(SB_T2_WEST_SB_OUT_B1_sel_inst0_O)
	);
	MuxWrapper_1_1 WIRE_SB_T0_EAST_SB_IN_B1(
		.I(SB_T0_EAST_SB_IN_B1),
		.O(WIRE_SB_T0_EAST_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T0_NORTH_SB_IN_B1(
		.I(SB_T0_NORTH_SB_IN_B1),
		.O(WIRE_SB_T0_NORTH_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T0_SOUTH_SB_IN_B1(
		.I(SB_T0_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T0_SOUTH_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T0_WEST_SB_IN_B1(
		.I(SB_T0_WEST_SB_IN_B1),
		.O(WIRE_SB_T0_WEST_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T1_EAST_SB_IN_B1(
		.I(SB_T1_EAST_SB_IN_B1),
		.O(WIRE_SB_T1_EAST_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T1_NORTH_SB_IN_B1(
		.I(SB_T1_NORTH_SB_IN_B1),
		.O(WIRE_SB_T1_NORTH_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T1_SOUTH_SB_IN_B1(
		.I(SB_T1_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T1_SOUTH_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T1_WEST_SB_IN_B1(
		.I(SB_T1_WEST_SB_IN_B1),
		.O(WIRE_SB_T1_WEST_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T2_EAST_SB_IN_B1(
		.I(SB_T2_EAST_SB_IN_B1),
		.O(WIRE_SB_T2_EAST_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T2_NORTH_SB_IN_B1(
		.I(SB_T2_NORTH_SB_IN_B1),
		.O(WIRE_SB_T2_NORTH_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T2_SOUTH_SB_IN_B1(
		.I(SB_T2_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T2_SOUTH_SB_IN_B1_O)
	);
	MuxWrapper_1_1 WIRE_SB_T2_WEST_SB_IN_B1(
		.I(SB_T2_WEST_SB_IN_B1),
		.O(WIRE_SB_T2_WEST_SB_IN_B1_O)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_18_32_inst0$bit_const_0_None(.out(ZextWrapper_18_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit18 ZextWrapper_18_32_inst0$self_I(
		.in(config_reg_1_O),
		.out(ZextWrapper_18_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_18_32_inst0$self_O_out;
	assign ZextWrapper_18_32_inst0$self_O_out = {ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$self_I_out[17:0]};
	mantle_wire__typeBitIn32 ZextWrapper_18_32_inst0$self_O(
		.in(ZextWrapper_18_32_inst0$self_O_in),
		.out(ZextWrapper_18_32_inst0$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_30_32_inst0$bit_const_0_None(.out(ZextWrapper_30_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit30 ZextWrapper_30_32_inst0$self_I(
		.in(config_reg_0_O),
		.out(ZextWrapper_30_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_30_32_inst0$self_O_out;
	assign ZextWrapper_30_32_inst0$self_O_out = {ZextWrapper_30_32_inst0$bit_const_0_None_out, ZextWrapper_30_32_inst0$bit_const_0_None_out, ZextWrapper_30_32_inst0$self_I_out[29:0]};
	mantle_wire__typeBitIn32 ZextWrapper_30_32_inst0$self_O(
		.in(ZextWrapper_30_32_inst0$self_O_in),
		.out(ZextWrapper_30_32_inst0$self_O_out)
	);
	coreir_and #(.width(1)) and1_inst0(
		.in0(coreir_eq_1_inst0_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst0_out)
	);
	coreir_and #(.width(1)) and1_inst1(
		.in0(coreir_eq_1_inst1_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst1_out)
	);
	coreir_and #(.width(1)) and1_inst10(
		.in0(coreir_eq_1_inst10_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst10_out)
	);
	coreir_and #(.width(1)) and1_inst11(
		.in0(coreir_eq_1_inst11_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst11_out)
	);
	coreir_and #(.width(1)) and1_inst2(
		.in0(coreir_eq_1_inst2_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst2_out)
	);
	coreir_and #(.width(1)) and1_inst3(
		.in0(coreir_eq_1_inst3_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst3_out)
	);
	coreir_and #(.width(1)) and1_inst4(
		.in0(coreir_eq_1_inst4_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst4_out)
	);
	coreir_and #(.width(1)) and1_inst5(
		.in0(coreir_eq_1_inst5_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst5_out)
	);
	coreir_and #(.width(1)) and1_inst6(
		.in0(coreir_eq_1_inst6_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst6_out)
	);
	coreir_and #(.width(1)) and1_inst7(
		.in0(coreir_eq_1_inst7_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst7_out)
	);
	coreir_and #(.width(1)) and1_inst8(
		.in0(coreir_eq_1_inst8_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst8_out)
	);
	coreir_and #(.width(1)) and1_inst9(
		.in0(coreir_eq_1_inst9_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst9_out)
	);
	ConfigRegister_30_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_18_8_32_1 config_reg_1(
		.clk(clk),
		.reset(reset),
		.O(config_reg_1_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	coreir_const #(
		.value(1'h1),
		.width(1)
	) const_1_1(.out(const_1_1_out));
	coreir_eq #(.width(1)) coreir_eq_1_inst0(
		.in0(const_1_1_out),
		.in1(RMUX_T0_NORTH_B1_sel_inst0_O),
		.out(coreir_eq_1_inst0_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst1(
		.in0(const_1_1_out),
		.in1(RMUX_T0_SOUTH_B1_sel_inst0_O),
		.out(coreir_eq_1_inst1_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst10(
		.in0(const_1_1_out),
		.in1(RMUX_T2_EAST_B1_sel_inst0_O),
		.out(coreir_eq_1_inst10_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst11(
		.in0(const_1_1_out),
		.in1(RMUX_T2_WEST_B1_sel_inst0_O),
		.out(coreir_eq_1_inst11_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst2(
		.in0(const_1_1_out),
		.in1(RMUX_T0_EAST_B1_sel_inst0_O),
		.out(coreir_eq_1_inst2_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst3(
		.in0(const_1_1_out),
		.in1(RMUX_T0_WEST_B1_sel_inst0_O),
		.out(coreir_eq_1_inst3_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst4(
		.in0(const_1_1_out),
		.in1(RMUX_T1_NORTH_B1_sel_inst0_O),
		.out(coreir_eq_1_inst4_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst5(
		.in0(const_1_1_out),
		.in1(RMUX_T1_SOUTH_B1_sel_inst0_O),
		.out(coreir_eq_1_inst5_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst6(
		.in0(const_1_1_out),
		.in1(RMUX_T1_EAST_B1_sel_inst0_O),
		.out(coreir_eq_1_inst6_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst7(
		.in0(const_1_1_out),
		.in1(RMUX_T1_WEST_B1_sel_inst0_O),
		.out(coreir_eq_1_inst7_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst8(
		.in0(const_1_1_out),
		.in1(RMUX_T2_NORTH_B1_sel_inst0_O),
		.out(coreir_eq_1_inst8_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst9(
		.in0(const_1_1_out),
		.in1(RMUX_T2_SOUTH_B1_sel_inst0_O),
		.out(coreir_eq_1_inst9_out)
	);
	assign SB_T0_EAST_SB_OUT_B1 = RMUX_T0_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T0_NORTH_SB_OUT_B1 = RMUX_T0_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T0_SOUTH_SB_OUT_B1 = RMUX_T0_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T0_WEST_SB_OUT_B1 = RMUX_T0_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T1_EAST_SB_OUT_B1 = RMUX_T1_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T1_NORTH_SB_OUT_B1 = RMUX_T1_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T1_SOUTH_SB_OUT_B1 = RMUX_T1_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T1_WEST_SB_OUT_B1 = RMUX_T1_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T2_EAST_SB_OUT_B1 = RMUX_T2_EAST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T2_NORTH_SB_OUT_B1 = RMUX_T2_NORTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T2_SOUTH_SB_OUT_B1 = RMUX_T2_SOUTH_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign SB_T2_WEST_SB_OUT_B1 = RMUX_T2_WEST_B1$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	assign read_config_data = MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
endmodule
module SB_ID0_3TRACKS_B16_MemCore (
	SB_T0_EAST_SB_IN_B16,
	SB_T0_EAST_SB_OUT_B16,
	SB_T0_NORTH_SB_IN_B16,
	SB_T0_NORTH_SB_OUT_B16,
	SB_T0_SOUTH_SB_IN_B16,
	SB_T0_SOUTH_SB_OUT_B16,
	SB_T0_WEST_SB_IN_B16,
	SB_T0_WEST_SB_OUT_B16,
	SB_T1_EAST_SB_IN_B16,
	SB_T1_EAST_SB_OUT_B16,
	SB_T1_NORTH_SB_IN_B16,
	SB_T1_NORTH_SB_OUT_B16,
	SB_T1_SOUTH_SB_IN_B16,
	SB_T1_SOUTH_SB_OUT_B16,
	SB_T1_WEST_SB_IN_B16,
	SB_T1_WEST_SB_OUT_B16,
	SB_T2_EAST_SB_IN_B16,
	SB_T2_EAST_SB_OUT_B16,
	SB_T2_NORTH_SB_IN_B16,
	SB_T2_NORTH_SB_OUT_B16,
	SB_T2_SOUTH_SB_IN_B16,
	SB_T2_SOUTH_SB_OUT_B16,
	SB_T2_WEST_SB_IN_B16,
	SB_T2_WEST_SB_OUT_B16,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	output_width_16_num_0,
	output_width_16_num_1,
	read_config_data,
	reset,
	stall
);
	input [15:0] SB_T0_EAST_SB_IN_B16;
	output [15:0] SB_T0_EAST_SB_OUT_B16;
	input [15:0] SB_T0_NORTH_SB_IN_B16;
	output [15:0] SB_T0_NORTH_SB_OUT_B16;
	input [15:0] SB_T0_SOUTH_SB_IN_B16;
	output [15:0] SB_T0_SOUTH_SB_OUT_B16;
	input [15:0] SB_T0_WEST_SB_IN_B16;
	output [15:0] SB_T0_WEST_SB_OUT_B16;
	input [15:0] SB_T1_EAST_SB_IN_B16;
	output [15:0] SB_T1_EAST_SB_OUT_B16;
	input [15:0] SB_T1_NORTH_SB_IN_B16;
	output [15:0] SB_T1_NORTH_SB_OUT_B16;
	input [15:0] SB_T1_SOUTH_SB_IN_B16;
	output [15:0] SB_T1_SOUTH_SB_OUT_B16;
	input [15:0] SB_T1_WEST_SB_IN_B16;
	output [15:0] SB_T1_WEST_SB_OUT_B16;
	input [15:0] SB_T2_EAST_SB_IN_B16;
	output [15:0] SB_T2_EAST_SB_OUT_B16;
	input [15:0] SB_T2_NORTH_SB_IN_B16;
	output [15:0] SB_T2_NORTH_SB_OUT_B16;
	input [15:0] SB_T2_SOUTH_SB_IN_B16;
	output [15:0] SB_T2_SOUTH_SB_OUT_B16;
	input [15:0] SB_T2_WEST_SB_IN_B16;
	output [15:0] SB_T2_WEST_SB_OUT_B16;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	input [15:0] output_width_16_num_0;
	input [15:0] output_width_16_num_1;
	output [31:0] read_config_data;
	input reset;
	input [0:0] stall;
	wire [0:0] Invert1_inst0_out;
	wire [15:0] MUX_SB_T0_EAST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out;
	wire [15:0] MUX_SB_T0_NORTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out;
	wire [15:0] MUX_SB_T0_SOUTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out;
	wire [15:0] MUX_SB_T0_WEST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out;
	wire [15:0] MUX_SB_T1_EAST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out;
	wire [15:0] MUX_SB_T1_NORTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out;
	wire [15:0] MUX_SB_T1_SOUTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out;
	wire [15:0] MUX_SB_T1_WEST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out;
	wire [15:0] MUX_SB_T2_EAST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out;
	wire [15:0] MUX_SB_T2_NORTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out;
	wire [15:0] MUX_SB_T2_SOUTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out;
	wire [15:0] MUX_SB_T2_WEST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out;
	wire [31:0] MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
	wire [15:0] REG_T0_EAST_B16_O;
	wire [15:0] REG_T0_NORTH_B16_O;
	wire [15:0] REG_T0_SOUTH_B16_O;
	wire [15:0] REG_T0_WEST_B16_O;
	wire [15:0] REG_T1_EAST_B16_O;
	wire [15:0] REG_T1_NORTH_B16_O;
	wire [15:0] REG_T1_SOUTH_B16_O;
	wire [15:0] REG_T1_WEST_B16_O;
	wire [15:0] REG_T2_EAST_B16_O;
	wire [15:0] REG_T2_NORTH_B16_O;
	wire [15:0] REG_T2_SOUTH_B16_O;
	wire [15:0] REG_T2_WEST_B16_O;
	wire [15:0] RMUX_T0_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T0_EAST_B16_sel_inst0_O;
	wire [15:0] RMUX_T0_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T0_NORTH_B16_sel_inst0_O;
	wire [15:0] RMUX_T0_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T0_SOUTH_B16_sel_inst0_O;
	wire [15:0] RMUX_T0_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T0_WEST_B16_sel_inst0_O;
	wire [15:0] RMUX_T1_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T1_EAST_B16_sel_inst0_O;
	wire [15:0] RMUX_T1_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T1_NORTH_B16_sel_inst0_O;
	wire [15:0] RMUX_T1_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T1_SOUTH_B16_sel_inst0_O;
	wire [15:0] RMUX_T1_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T1_WEST_B16_sel_inst0_O;
	wire [15:0] RMUX_T2_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T2_EAST_B16_sel_inst0_O;
	wire [15:0] RMUX_T2_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T2_NORTH_B16_sel_inst0_O;
	wire [15:0] RMUX_T2_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T2_SOUTH_B16_sel_inst0_O;
	wire [15:0] RMUX_T2_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [0:0] RMUX_T2_WEST_B16_sel_inst0_O;
	wire [2:0] SB_T0_EAST_SB_OUT_B16_sel_inst0_O;
	wire [2:0] SB_T0_NORTH_SB_OUT_B16_sel_inst0_O;
	wire [2:0] SB_T0_SOUTH_SB_OUT_B16_sel_inst0_O;
	wire [2:0] SB_T0_WEST_SB_OUT_B16_sel_inst0_O;
	wire [2:0] SB_T1_EAST_SB_OUT_B16_sel_inst0_O;
	wire [2:0] SB_T1_NORTH_SB_OUT_B16_sel_inst0_O;
	wire [2:0] SB_T1_SOUTH_SB_OUT_B16_sel_inst0_O;
	wire [2:0] SB_T1_WEST_SB_OUT_B16_sel_inst0_O;
	wire [2:0] SB_T2_EAST_SB_OUT_B16_sel_inst0_O;
	wire [2:0] SB_T2_NORTH_SB_OUT_B16_sel_inst0_O;
	wire [2:0] SB_T2_SOUTH_SB_OUT_B16_sel_inst0_O;
	wire [2:0] SB_T2_WEST_SB_OUT_B16_sel_inst0_O;
	wire [15:0] WIRE_SB_T0_EAST_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T0_NORTH_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T0_SOUTH_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T0_WEST_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T1_EAST_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T1_NORTH_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T1_SOUTH_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T1_WEST_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T2_EAST_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T2_NORTH_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T2_SOUTH_SB_IN_B16_O;
	wire [15:0] WIRE_SB_T2_WEST_SB_IN_B16_O;
	wire ZextWrapper_18_32_inst0$bit_const_0_None_out;
	wire [17:0] ZextWrapper_18_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_18_32_inst0$self_O_in;
	wire ZextWrapper_30_32_inst0$bit_const_0_None_out;
	wire [29:0] ZextWrapper_30_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_30_32_inst0$self_O_in;
	wire [0:0] and1_inst0_out;
	wire [0:0] and1_inst1_out;
	wire [0:0] and1_inst10_out;
	wire [0:0] and1_inst11_out;
	wire [0:0] and1_inst2_out;
	wire [0:0] and1_inst3_out;
	wire [0:0] and1_inst4_out;
	wire [0:0] and1_inst5_out;
	wire [0:0] and1_inst6_out;
	wire [0:0] and1_inst7_out;
	wire [0:0] and1_inst8_out;
	wire [0:0] and1_inst9_out;
	wire [29:0] config_reg_0_O;
	wire [17:0] config_reg_1_O;
	wire [0:0] const_1_1_out;
	wire coreir_eq_1_inst0_out;
	wire coreir_eq_1_inst1_out;
	wire coreir_eq_1_inst10_out;
	wire coreir_eq_1_inst11_out;
	wire coreir_eq_1_inst2_out;
	wire coreir_eq_1_inst3_out;
	wire coreir_eq_1_inst4_out;
	wire coreir_eq_1_inst5_out;
	wire coreir_eq_1_inst6_out;
	wire coreir_eq_1_inst7_out;
	wire coreir_eq_1_inst8_out;
	wire coreir_eq_1_inst9_out;
	coreir_not #(.width(1)) Invert1_inst0(
		.in(stall),
		.out(Invert1_inst0_out)
	);
	commonlib_muxn__N5__width16 MUX_SB_T0_EAST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0(
		.in_data_0(WIRE_SB_T0_WEST_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T2_NORTH_SB_IN_B16_O),
		.in_data_3(output_width_16_num_0),
		.in_data_4(output_width_16_num_1),
		.in_sel(SB_T0_EAST_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T0_EAST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out)
	);
	commonlib_muxn__N5__width16 MUX_SB_T0_NORTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0(
		.in_data_0(WIRE_SB_T0_WEST_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T1_EAST_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
		.in_data_3(output_width_16_num_0),
		.in_data_4(output_width_16_num_1),
		.in_sel(SB_T0_NORTH_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T0_NORTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out)
	);
	commonlib_muxn__N5__width16 MUX_SB_T0_SOUTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0(
		.in_data_0(WIRE_SB_T1_EAST_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T0_NORTH_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T1_WEST_SB_IN_B16_O),
		.in_data_3(output_width_16_num_0),
		.in_data_4(output_width_16_num_1),
		.in_sel(SB_T0_SOUTH_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T0_SOUTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out)
	);
	commonlib_muxn__N5__width16 MUX_SB_T0_WEST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0(
		.in_data_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
		.in_data_3(output_width_16_num_0),
		.in_data_4(output_width_16_num_1),
		.in_sel(SB_T0_WEST_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T0_WEST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out)
	);
	commonlib_muxn__N5__width16 MUX_SB_T1_EAST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0(
		.in_data_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T1_WEST_SB_IN_B16_O),
		.in_data_3(output_width_16_num_0),
		.in_data_4(output_width_16_num_1),
		.in_sel(SB_T1_EAST_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T1_EAST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out)
	);
	commonlib_muxn__N5__width16 MUX_SB_T1_NORTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0(
		.in_data_0(WIRE_SB_T2_EAST_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T2_WEST_SB_IN_B16_O),
		.in_data_3(output_width_16_num_0),
		.in_data_4(output_width_16_num_1),
		.in_sel(SB_T1_NORTH_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T1_NORTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out)
	);
	commonlib_muxn__N5__width16 MUX_SB_T1_SOUTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0(
		.in_data_0(WIRE_SB_T0_EAST_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T1_NORTH_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T2_WEST_SB_IN_B16_O),
		.in_data_3(output_width_16_num_0),
		.in_data_4(output_width_16_num_1),
		.in_sel(SB_T1_SOUTH_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T1_SOUTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out)
	);
	commonlib_muxn__N5__width16 MUX_SB_T1_WEST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0(
		.in_data_0(WIRE_SB_T2_NORTH_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T1_EAST_SB_IN_B16_O),
		.in_data_3(output_width_16_num_0),
		.in_data_4(output_width_16_num_1),
		.in_sel(SB_T1_WEST_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T1_WEST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out)
	);
	commonlib_muxn__N5__width16 MUX_SB_T2_EAST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0(
		.in_data_0(WIRE_SB_T1_NORTH_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T2_WEST_SB_IN_B16_O),
		.in_data_3(output_width_16_num_0),
		.in_data_4(output_width_16_num_1),
		.in_sel(SB_T2_EAST_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T2_EAST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out)
	);
	commonlib_muxn__N5__width16 MUX_SB_T2_NORTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0(
		.in_data_0(WIRE_SB_T1_WEST_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T0_EAST_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
		.in_data_3(output_width_16_num_0),
		.in_data_4(output_width_16_num_1),
		.in_sel(SB_T2_NORTH_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T2_NORTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out)
	);
	commonlib_muxn__N5__width16 MUX_SB_T2_SOUTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0(
		.in_data_0(WIRE_SB_T0_WEST_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T2_EAST_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T2_NORTH_SB_IN_B16_O),
		.in_data_3(output_width_16_num_0),
		.in_data_4(output_width_16_num_1),
		.in_sel(SB_T2_SOUTH_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T2_SOUTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out)
	);
	commonlib_muxn__N5__width16 MUX_SB_T2_WEST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0(
		.in_data_0(WIRE_SB_T1_NORTH_SB_IN_B16_O),
		.in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
		.in_data_2(WIRE_SB_T2_EAST_SB_IN_B16_O),
		.in_data_3(output_width_16_num_0),
		.in_data_4(output_width_16_num_1),
		.in_sel(SB_T2_WEST_SB_OUT_B16_sel_inst0_O),
		.out(MUX_SB_T2_WEST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out)
	);
	coreir_mux #(.width(32)) MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join(
		.in0(ZextWrapper_30_32_inst0$self_O_in),
		.in1(ZextWrapper_18_32_inst0$self_O_in),
		.sel(config_config_addr[0]),
		.out(MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out)
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_EAST_B16(
		.I(MUX_SB_T0_EAST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.O(REG_T0_EAST_B16_O),
		.CLK(clk),
		.CE(and1_inst2_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_NORTH_B16(
		.I(MUX_SB_T0_NORTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.O(REG_T0_NORTH_B16_O),
		.CLK(clk),
		.CE(and1_inst0_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_SOUTH_B16(
		.I(MUX_SB_T0_SOUTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.O(REG_T0_SOUTH_B16_O),
		.CLK(clk),
		.CE(and1_inst1_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_WEST_B16(
		.I(MUX_SB_T0_WEST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.O(REG_T0_WEST_B16_O),
		.CLK(clk),
		.CE(and1_inst3_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_EAST_B16(
		.I(MUX_SB_T1_EAST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.O(REG_T1_EAST_B16_O),
		.CLK(clk),
		.CE(and1_inst6_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_NORTH_B16(
		.I(MUX_SB_T1_NORTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.O(REG_T1_NORTH_B16_O),
		.CLK(clk),
		.CE(and1_inst4_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_SOUTH_B16(
		.I(MUX_SB_T1_SOUTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.O(REG_T1_SOUTH_B16_O),
		.CLK(clk),
		.CE(and1_inst5_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_WEST_B16(
		.I(MUX_SB_T1_WEST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.O(REG_T1_WEST_B16_O),
		.CLK(clk),
		.CE(and1_inst7_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_EAST_B16(
		.I(MUX_SB_T2_EAST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.O(REG_T2_EAST_B16_O),
		.CLK(clk),
		.CE(and1_inst10_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_NORTH_B16(
		.I(MUX_SB_T2_NORTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.O(REG_T2_NORTH_B16_O),
		.CLK(clk),
		.CE(and1_inst8_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_SOUTH_B16(
		.I(MUX_SB_T2_SOUTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.O(REG_T2_SOUTH_B16_O),
		.CLK(clk),
		.CE(and1_inst9_out[0])
	);
	Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_WEST_B16(
		.I(MUX_SB_T2_WEST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.O(REG_T2_WEST_B16_O),
		.CLK(clk),
		.CE(and1_inst11_out[0])
	);
	coreir_mux #(.width(16)) RMUX_T0_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T0_EAST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.in1(REG_T0_EAST_B16_O),
		.sel(RMUX_T0_EAST_B16_sel_inst0_O[0]),
		.out(RMUX_T0_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T0_EAST_B16_sel_unq1 RMUX_T0_EAST_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T0_EAST_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T0_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T0_NORTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.in1(REG_T0_NORTH_B16_O),
		.sel(RMUX_T0_NORTH_B16_sel_inst0_O[0]),
		.out(RMUX_T0_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T0_NORTH_B16_sel_unq1 RMUX_T0_NORTH_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T0_NORTH_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T0_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T0_SOUTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.in1(REG_T0_SOUTH_B16_O),
		.sel(RMUX_T0_SOUTH_B16_sel_inst0_O[0]),
		.out(RMUX_T0_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T0_SOUTH_B16_sel_unq1 RMUX_T0_SOUTH_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T0_SOUTH_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T0_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T0_WEST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.in1(REG_T0_WEST_B16_O),
		.sel(RMUX_T0_WEST_B16_sel_inst0_O[0]),
		.out(RMUX_T0_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T0_WEST_B16_sel_unq1 RMUX_T0_WEST_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T0_WEST_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T1_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T1_EAST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.in1(REG_T1_EAST_B16_O),
		.sel(RMUX_T1_EAST_B16_sel_inst0_O[0]),
		.out(RMUX_T1_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T1_EAST_B16_sel_unq1 RMUX_T1_EAST_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T1_EAST_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T1_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T1_NORTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.in1(REG_T1_NORTH_B16_O),
		.sel(RMUX_T1_NORTH_B16_sel_inst0_O[0]),
		.out(RMUX_T1_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T1_NORTH_B16_sel_unq1 RMUX_T1_NORTH_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T1_NORTH_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T1_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T1_SOUTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.in1(REG_T1_SOUTH_B16_O),
		.sel(RMUX_T1_SOUTH_B16_sel_inst0_O[0]),
		.out(RMUX_T1_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T1_SOUTH_B16_sel_unq1 RMUX_T1_SOUTH_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T1_SOUTH_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T1_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T1_WEST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.in1(REG_T1_WEST_B16_O),
		.sel(RMUX_T1_WEST_B16_sel_inst0_O[0]),
		.out(RMUX_T1_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T1_WEST_B16_sel_unq1 RMUX_T1_WEST_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T1_WEST_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T2_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T2_EAST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.in1(REG_T2_EAST_B16_O),
		.sel(RMUX_T2_EAST_B16_sel_inst0_O[0]),
		.out(RMUX_T2_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T2_EAST_B16_sel_unq1 RMUX_T2_EAST_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T2_EAST_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T2_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T2_NORTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.in1(REG_T2_NORTH_B16_O),
		.sel(RMUX_T2_NORTH_B16_sel_inst0_O[0]),
		.out(RMUX_T2_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T2_NORTH_B16_sel_unq1 RMUX_T2_NORTH_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T2_NORTH_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T2_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T2_SOUTH_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.in1(REG_T2_SOUTH_B16_O),
		.sel(RMUX_T2_SOUTH_B16_sel_inst0_O[0]),
		.out(RMUX_T2_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T2_SOUTH_B16_sel_unq1 RMUX_T2_SOUTH_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T2_SOUTH_B16_sel_inst0_O)
	);
	coreir_mux #(.width(16)) RMUX_T2_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(MUX_SB_T2_WEST_SB_OUT_B16$Mux5xBits16_inst0$coreir_commonlib_mux5x16_inst0_out),
		.in1(REG_T2_WEST_B16_O),
		.sel(RMUX_T2_WEST_B16_sel_inst0_O[0]),
		.out(RMUX_T2_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	RMUX_T2_WEST_B16_sel_unq1 RMUX_T2_WEST_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(RMUX_T2_WEST_B16_sel_inst0_O)
	);
	SB_T0_EAST_SB_OUT_B16_sel_unq1 SB_T0_EAST_SB_OUT_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T0_EAST_SB_OUT_B16_sel_inst0_O)
	);
	SB_T0_NORTH_SB_OUT_B16_sel_unq1 SB_T0_NORTH_SB_OUT_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T0_NORTH_SB_OUT_B16_sel_inst0_O)
	);
	SB_T0_SOUTH_SB_OUT_B16_sel_unq1 SB_T0_SOUTH_SB_OUT_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T0_SOUTH_SB_OUT_B16_sel_inst0_O)
	);
	SB_T0_WEST_SB_OUT_B16_sel_unq1 SB_T0_WEST_SB_OUT_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T0_WEST_SB_OUT_B16_sel_inst0_O)
	);
	SB_T1_EAST_SB_OUT_B16_sel_unq1 SB_T1_EAST_SB_OUT_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T1_EAST_SB_OUT_B16_sel_inst0_O)
	);
	SB_T1_NORTH_SB_OUT_B16_sel_unq1 SB_T1_NORTH_SB_OUT_B16_sel_inst0(
		.I(config_reg_0_O),
		.O(SB_T1_NORTH_SB_OUT_B16_sel_inst0_O)
	);
	SB_T1_SOUTH_SB_OUT_B16_sel_unq1 SB_T1_SOUTH_SB_OUT_B16_sel_inst0(
		.I(config_reg_1_O),
		.O(SB_T1_SOUTH_SB_OUT_B16_sel_inst0_O)
	);
	SB_T1_WEST_SB_OUT_B16_sel_unq1 SB_T1_WEST_SB_OUT_B16_sel_inst0(
		.I(config_reg_1_O),
		.O(SB_T1_WEST_SB_OUT_B16_sel_inst0_O)
	);
	SB_T2_EAST_SB_OUT_B16_sel_unq1 SB_T2_EAST_SB_OUT_B16_sel_inst0(
		.I(config_reg_1_O),
		.O(SB_T2_EAST_SB_OUT_B16_sel_inst0_O)
	);
	SB_T2_NORTH_SB_OUT_B16_sel_unq1 SB_T2_NORTH_SB_OUT_B16_sel_inst0(
		.I(config_reg_1_O),
		.O(SB_T2_NORTH_SB_OUT_B16_sel_inst0_O)
	);
	SB_T2_SOUTH_SB_OUT_B16_sel_unq1 SB_T2_SOUTH_SB_OUT_B16_sel_inst0(
		.I(config_reg_1_O),
		.O(SB_T2_SOUTH_SB_OUT_B16_sel_inst0_O)
	);
	SB_T2_WEST_SB_OUT_B16_sel_unq1 SB_T2_WEST_SB_OUT_B16_sel_inst0(
		.I(config_reg_1_O),
		.O(SB_T2_WEST_SB_OUT_B16_sel_inst0_O)
	);
	MuxWrapper_1_16 WIRE_SB_T0_EAST_SB_IN_B16(
		.I(SB_T0_EAST_SB_IN_B16),
		.O(WIRE_SB_T0_EAST_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T0_NORTH_SB_IN_B16(
		.I(SB_T0_NORTH_SB_IN_B16),
		.O(WIRE_SB_T0_NORTH_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T0_SOUTH_SB_IN_B16(
		.I(SB_T0_SOUTH_SB_IN_B16),
		.O(WIRE_SB_T0_SOUTH_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T0_WEST_SB_IN_B16(
		.I(SB_T0_WEST_SB_IN_B16),
		.O(WIRE_SB_T0_WEST_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T1_EAST_SB_IN_B16(
		.I(SB_T1_EAST_SB_IN_B16),
		.O(WIRE_SB_T1_EAST_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T1_NORTH_SB_IN_B16(
		.I(SB_T1_NORTH_SB_IN_B16),
		.O(WIRE_SB_T1_NORTH_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T1_SOUTH_SB_IN_B16(
		.I(SB_T1_SOUTH_SB_IN_B16),
		.O(WIRE_SB_T1_SOUTH_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T1_WEST_SB_IN_B16(
		.I(SB_T1_WEST_SB_IN_B16),
		.O(WIRE_SB_T1_WEST_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T2_EAST_SB_IN_B16(
		.I(SB_T2_EAST_SB_IN_B16),
		.O(WIRE_SB_T2_EAST_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T2_NORTH_SB_IN_B16(
		.I(SB_T2_NORTH_SB_IN_B16),
		.O(WIRE_SB_T2_NORTH_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T2_SOUTH_SB_IN_B16(
		.I(SB_T2_SOUTH_SB_IN_B16),
		.O(WIRE_SB_T2_SOUTH_SB_IN_B16_O)
	);
	MuxWrapper_1_16 WIRE_SB_T2_WEST_SB_IN_B16(
		.I(SB_T2_WEST_SB_IN_B16),
		.O(WIRE_SB_T2_WEST_SB_IN_B16_O)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_18_32_inst0$bit_const_0_None(.out(ZextWrapper_18_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit18 ZextWrapper_18_32_inst0$self_I(
		.in(config_reg_1_O),
		.out(ZextWrapper_18_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_18_32_inst0$self_O_out;
	assign ZextWrapper_18_32_inst0$self_O_out = {ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$bit_const_0_None_out, ZextWrapper_18_32_inst0$self_I_out[17:0]};
	mantle_wire__typeBitIn32 ZextWrapper_18_32_inst0$self_O(
		.in(ZextWrapper_18_32_inst0$self_O_in),
		.out(ZextWrapper_18_32_inst0$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_30_32_inst0$bit_const_0_None(.out(ZextWrapper_30_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit30 ZextWrapper_30_32_inst0$self_I(
		.in(config_reg_0_O),
		.out(ZextWrapper_30_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_30_32_inst0$self_O_out;
	assign ZextWrapper_30_32_inst0$self_O_out = {ZextWrapper_30_32_inst0$bit_const_0_None_out, ZextWrapper_30_32_inst0$bit_const_0_None_out, ZextWrapper_30_32_inst0$self_I_out[29:0]};
	mantle_wire__typeBitIn32 ZextWrapper_30_32_inst0$self_O(
		.in(ZextWrapper_30_32_inst0$self_O_in),
		.out(ZextWrapper_30_32_inst0$self_O_out)
	);
	coreir_and #(.width(1)) and1_inst0(
		.in0(coreir_eq_1_inst0_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst0_out)
	);
	coreir_and #(.width(1)) and1_inst1(
		.in0(coreir_eq_1_inst1_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst1_out)
	);
	coreir_and #(.width(1)) and1_inst10(
		.in0(coreir_eq_1_inst10_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst10_out)
	);
	coreir_and #(.width(1)) and1_inst11(
		.in0(coreir_eq_1_inst11_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst11_out)
	);
	coreir_and #(.width(1)) and1_inst2(
		.in0(coreir_eq_1_inst2_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst2_out)
	);
	coreir_and #(.width(1)) and1_inst3(
		.in0(coreir_eq_1_inst3_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst3_out)
	);
	coreir_and #(.width(1)) and1_inst4(
		.in0(coreir_eq_1_inst4_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst4_out)
	);
	coreir_and #(.width(1)) and1_inst5(
		.in0(coreir_eq_1_inst5_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst5_out)
	);
	coreir_and #(.width(1)) and1_inst6(
		.in0(coreir_eq_1_inst6_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst6_out)
	);
	coreir_and #(.width(1)) and1_inst7(
		.in0(coreir_eq_1_inst7_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst7_out)
	);
	coreir_and #(.width(1)) and1_inst8(
		.in0(coreir_eq_1_inst8_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst8_out)
	);
	coreir_and #(.width(1)) and1_inst9(
		.in0(coreir_eq_1_inst9_out),
		.in1(Invert1_inst0_out),
		.out(and1_inst9_out)
	);
	ConfigRegister_30_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_18_8_32_1 config_reg_1(
		.clk(clk),
		.reset(reset),
		.O(config_reg_1_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	coreir_const #(
		.value(1'h1),
		.width(1)
	) const_1_1(.out(const_1_1_out));
	coreir_eq #(.width(1)) coreir_eq_1_inst0(
		.in0(const_1_1_out),
		.in1(RMUX_T0_NORTH_B16_sel_inst0_O),
		.out(coreir_eq_1_inst0_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst1(
		.in0(const_1_1_out),
		.in1(RMUX_T0_SOUTH_B16_sel_inst0_O),
		.out(coreir_eq_1_inst1_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst10(
		.in0(const_1_1_out),
		.in1(RMUX_T2_EAST_B16_sel_inst0_O),
		.out(coreir_eq_1_inst10_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst11(
		.in0(const_1_1_out),
		.in1(RMUX_T2_WEST_B16_sel_inst0_O),
		.out(coreir_eq_1_inst11_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst2(
		.in0(const_1_1_out),
		.in1(RMUX_T0_EAST_B16_sel_inst0_O),
		.out(coreir_eq_1_inst2_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst3(
		.in0(const_1_1_out),
		.in1(RMUX_T0_WEST_B16_sel_inst0_O),
		.out(coreir_eq_1_inst3_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst4(
		.in0(const_1_1_out),
		.in1(RMUX_T1_NORTH_B16_sel_inst0_O),
		.out(coreir_eq_1_inst4_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst5(
		.in0(const_1_1_out),
		.in1(RMUX_T1_SOUTH_B16_sel_inst0_O),
		.out(coreir_eq_1_inst5_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst6(
		.in0(const_1_1_out),
		.in1(RMUX_T1_EAST_B16_sel_inst0_O),
		.out(coreir_eq_1_inst6_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst7(
		.in0(const_1_1_out),
		.in1(RMUX_T1_WEST_B16_sel_inst0_O),
		.out(coreir_eq_1_inst7_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst8(
		.in0(const_1_1_out),
		.in1(RMUX_T2_NORTH_B16_sel_inst0_O),
		.out(coreir_eq_1_inst8_out)
	);
	coreir_eq #(.width(1)) coreir_eq_1_inst9(
		.in0(const_1_1_out),
		.in1(RMUX_T2_SOUTH_B16_sel_inst0_O),
		.out(coreir_eq_1_inst9_out)
	);
	assign SB_T0_EAST_SB_OUT_B16 = RMUX_T0_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T0_NORTH_SB_OUT_B16 = RMUX_T0_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T0_SOUTH_SB_OUT_B16 = RMUX_T0_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T0_WEST_SB_OUT_B16 = RMUX_T0_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T1_EAST_SB_OUT_B16 = RMUX_T1_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T1_NORTH_SB_OUT_B16 = RMUX_T1_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T1_SOUTH_SB_OUT_B16 = RMUX_T1_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T1_WEST_SB_OUT_B16 = RMUX_T1_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T2_EAST_SB_OUT_B16 = RMUX_T2_EAST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T2_NORTH_SB_OUT_B16 = RMUX_T2_NORTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T2_SOUTH_SB_OUT_B16 = RMUX_T2_SOUTH_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign SB_T2_WEST_SB_OUT_B16 = RMUX_T2_WEST_B16$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	assign read_config_data = MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
endmodule
module ConfigRegister_17_8_32_75 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [16:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [16:0] Register_inst0_O;
	wire [7:0] const_75_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq5 Register_inst0(
		.I(config_data[16:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h4b),
		.width(8)
	) const_75_8(.out(const_75_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_75_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_17_8_32_59 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [16:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [16:0] Register_inst0_O;
	wire [7:0] const_59_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq5 Register_inst0(
		.I(config_data[16:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h3b),
		.width(8)
	) const_59_8(.out(const_59_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_59_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_17_8_32_55 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [16:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [16:0] Register_inst0_O;
	wire [7:0] const_55_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq5 Register_inst0(
		.I(config_data[16:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h37),
		.width(8)
	) const_55_8(.out(const_55_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_55_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_17_8_32_30 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [16:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [16:0] Register_inst0_O;
	wire [7:0] const_30_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq5 Register_inst0(
		.I(config_data[16:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h1e),
		.width(8)
	) const_30_8(.out(const_30_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_30_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_17_8_32_3 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [16:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [16:0] Register_inst0_O;
	wire [7:0] const_3_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq5 Register_inst0(
		.I(config_data[16:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h03),
		.width(8)
	) const_3_8(.out(const_3_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_3_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_17_8_32_26 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [16:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [16:0] Register_inst0_O;
	wire [7:0] const_26_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq5 Register_inst0(
		.I(config_data[16:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h1a),
		.width(8)
	) const_26_8(.out(const_26_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_26_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_17_8_32_15 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [16:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [16:0] Register_inst0_O;
	wire [7:0] const_15_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq5 Register_inst0(
		.I(config_data[16:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h0f),
		.width(8)
	) const_15_8(.out(const_15_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_15_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_17_8_32_11 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [16:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [16:0] Register_inst0_O;
	wire [7:0] const_11_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq5 Register_inst0(
		.I(config_data[16:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h0b),
		.width(8)
	) const_11_8(.out(const_11_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_11_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module ConfigRegister_11_8_32_81 (
	clk,
	reset,
	O,
	config_addr,
	config_data,
	config_en
);
	input clk;
	input reset;
	output [10:0] O;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	wire [10:0] Register_inst0_O;
	wire [7:0] const_81_8_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bits_8_eq_inst0_out;
	Register_unq9 Register_inst0(
		.I(config_data[10:0]),
		.O(Register_inst0_O),
		.CE(magma_Bit_and_inst0_out),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	coreir_const #(
		.value(8'h51),
		.width(8)
	) const_81_8(.out(const_81_8_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(config_addr),
		.in1(const_81_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	assign O = Register_inst0_O;
endmodule
module MemCore (
	clk,
	config_1_config_addr,
	config_1_config_data,
	config_1_read,
	config_1_write,
	config_config_addr,
	config_config_data,
	config_en_0,
	config_read,
	config_write,
	flush,
	input_width_16_num_0,
	input_width_16_num_1,
	input_width_16_num_2,
	input_width_16_num_3,
	input_width_1_num_0,
	input_width_1_num_1,
	output_width_16_num_0,
	output_width_16_num_1,
	output_width_1_num_0,
	output_width_1_num_1,
	output_width_1_num_2,
	read_config_data,
	read_config_data_1,
	reset,
	stall
);
	input clk;
	input [7:0] config_1_config_addr;
	input [31:0] config_1_config_data;
	input [0:0] config_1_read;
	input [0:0] config_1_write;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input config_en_0;
	input [0:0] config_read;
	input [0:0] config_write;
	input [0:0] flush;
	input [15:0] input_width_16_num_0;
	input [15:0] input_width_16_num_1;
	input [15:0] input_width_16_num_2;
	input [15:0] input_width_16_num_3;
	input [0:0] input_width_1_num_0;
	input [0:0] input_width_1_num_1;
	output [15:0] output_width_16_num_0;
	output [15:0] output_width_16_num_1;
	output [0:0] output_width_1_num_0;
	output [0:0] output_width_1_num_1;
	output [0:0] output_width_1_num_2;
	output [31:0] read_config_data;
	output [31:0] read_config_data_1;
	input reset;
	input [0:0] stall;
	wire [0:0] AND_CONFIG_EN_SRAM_0_out;
	wire [0:0] Invert1_inst0_out;
	wire [0:0] Invert1_inst1_out;
	wire [0:0] LakeTop_W_inst0_output_width_1_num_1;
	wire [0:0] LakeTop_W_inst0_output_width_1_num_0;
	wire [15:0] LakeTop_W_inst0_output_width_16_num_1;
	wire [15:0] LakeTop_W_inst0_output_width_16_num_0;
	wire [0:0] LakeTop_W_inst0_output_width_1_num_2;
	wire [31:0] LakeTop_W_inst0_config_data_out;
	wire [31:0] MuxWrapper_82_32_inst0$Mux82xBits32_inst0$coreir_commonlib_mux82x32_inst0_out;
	wire [6:0] MuxWrapper_82_32_inst0_S_in;
	wire [0:0] OR_CONFIG_EN_SRAM_0_out;
	wire OR_CONFIG_RD_SRAM$orr_inst0_out;
	wire OR_CONFIG_WR_SRAM$orr_inst0_out;
	wire [7:0] OR_config_addr_FEATURE_out;
	wire [31:0] OR_config_data_FEATURE_out;
	wire ZextWrapper_11_32_inst0$bit_const_0_None_out;
	wire [10:0] ZextWrapper_11_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_11_32_inst0$self_O_in;
	wire ZextWrapper_17_32_inst0$bit_const_0_None_out;
	wire [16:0] ZextWrapper_17_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_17_32_inst0$self_O_in;
	wire ZextWrapper_17_32_inst1$bit_const_0_None_out;
	wire [16:0] ZextWrapper_17_32_inst1$self_I_out;
	wire [31:0] ZextWrapper_17_32_inst1$self_O_in;
	wire ZextWrapper_17_32_inst2$bit_const_0_None_out;
	wire [16:0] ZextWrapper_17_32_inst2$self_I_out;
	wire [31:0] ZextWrapper_17_32_inst2$self_O_in;
	wire ZextWrapper_17_32_inst3$bit_const_0_None_out;
	wire [16:0] ZextWrapper_17_32_inst3$self_I_out;
	wire [31:0] ZextWrapper_17_32_inst3$self_O_in;
	wire ZextWrapper_17_32_inst4$bit_const_0_None_out;
	wire [16:0] ZextWrapper_17_32_inst4$self_I_out;
	wire [31:0] ZextWrapper_17_32_inst4$self_O_in;
	wire ZextWrapper_17_32_inst5$bit_const_0_None_out;
	wire [16:0] ZextWrapper_17_32_inst5$self_I_out;
	wire [31:0] ZextWrapper_17_32_inst5$self_O_in;
	wire ZextWrapper_17_32_inst6$bit_const_0_None_out;
	wire [16:0] ZextWrapper_17_32_inst6$self_I_out;
	wire [31:0] ZextWrapper_17_32_inst6$self_O_in;
	wire ZextWrapper_17_32_inst7$bit_const_0_None_out;
	wire [16:0] ZextWrapper_17_32_inst7$self_I_out;
	wire [31:0] ZextWrapper_17_32_inst7$self_O_in;
	wire ZextWrapper_20_32_inst0$bit_const_0_None_out;
	wire [19:0] ZextWrapper_20_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_20_32_inst0$self_O_in;
	wire ZextWrapper_20_32_inst1$bit_const_0_None_out;
	wire [19:0] ZextWrapper_20_32_inst1$self_I_out;
	wire [31:0] ZextWrapper_20_32_inst1$self_O_in;
	wire ZextWrapper_20_32_inst2$bit_const_0_None_out;
	wire [19:0] ZextWrapper_20_32_inst2$self_I_out;
	wire [31:0] ZextWrapper_20_32_inst2$self_O_in;
	wire ZextWrapper_20_32_inst3$bit_const_0_None_out;
	wire [19:0] ZextWrapper_20_32_inst3$self_I_out;
	wire [31:0] ZextWrapper_20_32_inst3$self_O_in;
	wire ZextWrapper_20_32_inst4$bit_const_0_None_out;
	wire [19:0] ZextWrapper_20_32_inst4$self_I_out;
	wire [31:0] ZextWrapper_20_32_inst4$self_O_in;
	wire ZextWrapper_20_32_inst5$bit_const_0_None_out;
	wire [19:0] ZextWrapper_20_32_inst5$self_I_out;
	wire [31:0] ZextWrapper_20_32_inst5$self_O_in;
	wire ZextWrapper_20_32_inst6$bit_const_0_None_out;
	wire [19:0] ZextWrapper_20_32_inst6$self_I_out;
	wire [31:0] ZextWrapper_20_32_inst6$self_O_in;
	wire ZextWrapper_25_32_inst0$bit_const_0_None_out;
	wire [24:0] ZextWrapper_25_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_25_32_inst0$self_O_in;
	wire ZextWrapper_25_32_inst1$bit_const_0_None_out;
	wire [24:0] ZextWrapper_25_32_inst1$self_I_out;
	wire [31:0] ZextWrapper_25_32_inst1$self_O_in;
	wire ZextWrapper_26_32_inst0$bit_const_0_None_out;
	wire [25:0] ZextWrapper_26_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_26_32_inst0$self_O_in;
	wire ZextWrapper_28_32_inst0$bit_const_0_None_out;
	wire [27:0] ZextWrapper_28_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_28_32_inst0$self_O_in;
	wire [25:0] config_reg_0_O;
	wire [31:0] config_reg_1_O;
	wire [31:0] config_reg_10_O;
	wire [16:0] config_reg_11_O;
	wire [31:0] config_reg_12_O;
	wire [31:0] config_reg_13_O;
	wire [31:0] config_reg_14_O;
	wire [16:0] config_reg_15_O;
	wire [31:0] config_reg_16_O;
	wire [31:0] config_reg_17_O;
	wire [31:0] config_reg_18_O;
	wire [19:0] config_reg_19_O;
	wire [31:0] config_reg_2_O;
	wire [31:0] config_reg_20_O;
	wire [31:0] config_reg_21_O;
	wire [19:0] config_reg_22_O;
	wire [31:0] config_reg_23_O;
	wire [31:0] config_reg_24_O;
	wire [31:0] config_reg_25_O;
	wire [16:0] config_reg_26_O;
	wire [31:0] config_reg_27_O;
	wire [31:0] config_reg_28_O;
	wire [31:0] config_reg_29_O;
	wire [16:0] config_reg_3_O;
	wire [16:0] config_reg_30_O;
	wire [31:0] config_reg_31_O;
	wire [31:0] config_reg_32_O;
	wire [31:0] config_reg_33_O;
	wire [19:0] config_reg_34_O;
	wire [31:0] config_reg_35_O;
	wire [31:0] config_reg_36_O;
	wire [19:0] config_reg_37_O;
	wire [31:0] config_reg_38_O;
	wire [31:0] config_reg_39_O;
	wire [31:0] config_reg_4_O;
	wire [31:0] config_reg_40_O;
	wire [24:0] config_reg_41_O;
	wire [31:0] config_reg_42_O;
	wire [31:0] config_reg_43_O;
	wire [31:0] config_reg_44_O;
	wire [31:0] config_reg_45_O;
	wire [31:0] config_reg_46_O;
	wire [31:0] config_reg_47_O;
	wire [27:0] config_reg_48_O;
	wire [31:0] config_reg_49_O;
	wire [31:0] config_reg_5_O;
	wire [31:0] config_reg_50_O;
	wire [19:0] config_reg_51_O;
	wire [31:0] config_reg_52_O;
	wire [31:0] config_reg_53_O;
	wire [31:0] config_reg_54_O;
	wire [16:0] config_reg_55_O;
	wire [31:0] config_reg_56_O;
	wire [31:0] config_reg_57_O;
	wire [31:0] config_reg_58_O;
	wire [16:0] config_reg_59_O;
	wire [31:0] config_reg_6_O;
	wire [31:0] config_reg_60_O;
	wire [31:0] config_reg_61_O;
	wire [31:0] config_reg_62_O;
	wire [19:0] config_reg_63_O;
	wire [31:0] config_reg_64_O;
	wire [31:0] config_reg_65_O;
	wire [19:0] config_reg_66_O;
	wire [31:0] config_reg_67_O;
	wire [31:0] config_reg_68_O;
	wire [31:0] config_reg_69_O;
	wire [31:0] config_reg_7_O;
	wire [31:0] config_reg_70_O;
	wire [24:0] config_reg_71_O;
	wire [31:0] config_reg_72_O;
	wire [31:0] config_reg_73_O;
	wire [31:0] config_reg_74_O;
	wire [16:0] config_reg_75_O;
	wire [31:0] config_reg_76_O;
	wire [31:0] config_reg_77_O;
	wire [31:0] config_reg_78_O;
	wire [31:0] config_reg_79_O;
	wire [31:0] config_reg_8_O;
	wire [31:0] config_reg_80_O;
	wire [10:0] config_reg_81_O;
	wire [31:0] config_reg_9_O;
	wire coreir_wrapInAsyncReset_inst0_out;
	wire coreir_wrapOutAsyncReset_inst0_out;
	wire [0:0] flush_reg_sel_inst0_O;
	wire [0:0] flush_reg_value_inst0_O;
	wire [0:0] flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] input_width_1_num_0_reg_sel_inst0_O;
	wire [0:0] input_width_1_num_0_reg_value_inst0_O;
	wire [0:0] input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] input_width_1_num_1_reg_sel_inst0_O;
	wire [0:0] input_width_1_num_1_reg_value_inst0_O;
	wire [0:0] input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [3:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality_inst0_O;
	wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0_inst0_O;
	wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1_inst0_O;
	wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2_inst0_O;
	wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3_inst0_O;
	wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4_inst0_O;
	wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5_inst0_O;
	wire [0:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable_inst0_O;
	wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr_inst0_O;
	wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0_inst0_O;
	wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1_inst0_O;
	wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2_inst0_O;
	wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3_inst0_O;
	wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4_inst0_O;
	wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_0_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_1_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_2_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_3_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_4_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_5_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_0_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_1_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_2_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_3_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_4_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_5_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_3_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_4_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_5_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_3_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_4_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_5_inst0_O;
	wire [0:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5_inst0_O;
	wire [0:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_3_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_4_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_5_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_3_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_4_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_5_inst0_O;
	wire [0:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5_inst0_O;
	wire [0:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5_inst0_O;
	wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4_inst0_O;
	wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5_inst0_O;
	wire [0:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_0_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_1_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_2_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_3_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_4_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_5_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_0_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_1_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_2_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_3_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_4_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_5_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4_inst0_O;
	wire [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5_inst0_O;
	// wire [0:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5_inst0_O;
	// wire [0:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5_inst0_O;
	// wire [0:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5_inst0_O;
	// wire [0:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4_inst0_O;
	// wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4_inst0_O;
	// wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5_inst0_O;
	wire [1:0] mode_inst0_O;
	wire [7:0] self_config_config_addr_out;
	wire [0:0] tile_en_inst0_O;
	coreir_and #(.width(1)) AND_CONFIG_EN_SRAM_0(
		.in0(OR_CONFIG_EN_SRAM_0_out),
		.in1(config_en_0),
		.out(AND_CONFIG_EN_SRAM_0_out)
	);
	coreir_not #(.width(1)) Invert1_inst0(
		.in(coreir_wrapInAsyncReset_inst0_out),
		.out(Invert1_inst0_out)
	);
	coreir_not #(.width(1)) Invert1_inst1(
		.in(stall),
		.out(Invert1_inst1_out)
	);
	LakeTop_W LakeTop_W_inst0(
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_0_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2_inst0_O),
		.mode(mode_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_5_inst0_O),
		.mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable_inst0_O),
		.input_width_16_num_3(input_width_16_num_3),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5_inst0_O),
		.mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5_inst0_O),
		.output_width_1_num_1(LakeTop_W_inst0_output_width_1_num_1),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_1_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en_inst0_O),
		.mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_4_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_3_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1_inst0_O),
		.output_width_1_num_0(LakeTop_W_inst0_output_width_1_num_0),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_1_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1_inst0_O),
		.mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_4_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2_inst0_O),
		.mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_1_inst0_O),
		.config_en(AND_CONFIG_EN_SRAM_0_out),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_0_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_2_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_3_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality_inst0_O),
		.output_width_16_num_1(LakeTop_W_inst0_output_width_16_num_1),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_2_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_5_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_3_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_3_inst0_O),
		.mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5_inst0_O),
		.input_width_16_num_0(input_width_16_num_0),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1_inst0_O),
		.config_write(OR_CONFIG_RD_SRAM$orr_inst0_out),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_3_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_5_inst0_O),
		.mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_3_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2_inst0_O),
		.clk(clk),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_0_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0_inst0_O),
		.mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0_inst0_O),
		.flush(flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality_inst0_O),
		.output_width_16_num_0(LakeTop_W_inst0_output_width_16_num_0),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1_inst0_O),
		.output_width_1_num_2(LakeTop_W_inst0_output_width_1_num_2),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_4_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_4_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0_inst0_O),
		.clk_en(Invert1_inst1_out),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable_inst0_O),
		.rst_n(coreir_wrapOutAsyncReset_inst0_out),
		.config_read(OR_CONFIG_WR_SRAM$orr_inst0_out),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2_inst0_O),
		.input_width_1_num_0(input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_5_inst0_O),
		.input_width_16_num_2(input_width_16_num_2),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4_inst0_O),
		.config_data_in(OR_config_data_FEATURE_out),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_4_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2_inst0_O),
		.mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5_inst0_O),
		.input_width_1_num_1(input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_4_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4_inst0_O),
		.tile_en(tile_en_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1_inst0_O),
		.mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_2_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_4_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_4_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_5_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_5_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0_inst0_O),
		.config_addr_in(OR_config_addr_FEATURE_out),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_1_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0_inst0_O),
		.mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_3_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable_inst0_O),
		.config_data_out(LakeTop_W_inst0_config_data_out),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_5_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5_inst0_O),
		.input_width_16_num_1(input_width_16_num_1),
		.mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3_inst0_O),
		.mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr_inst0_O),
		// .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_2_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_0_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_3_inst0_O),
		.mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_5_inst0_O),
		.mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1_inst0_O)
	);
	commonlib_muxn__N82__width32 MuxWrapper_82_32_inst0$Mux82xBits32_inst0$coreir_commonlib_mux82x32_inst0(
		.in_data_0(ZextWrapper_26_32_inst0$self_O_in),
		.in_data_1(config_reg_1_O),
		.in_data_10(config_reg_10_O),
		.in_data_11(ZextWrapper_17_32_inst1$self_O_in),
		.in_data_12(config_reg_12_O),
		.in_data_13(config_reg_13_O),
		.in_data_14(config_reg_14_O),
		.in_data_15(ZextWrapper_17_32_inst2$self_O_in),
		.in_data_16(config_reg_16_O),
		.in_data_17(config_reg_17_O),
		.in_data_18(config_reg_18_O),
		.in_data_19(ZextWrapper_20_32_inst0$self_O_in),
		.in_data_2(config_reg_2_O),
		.in_data_20(config_reg_20_O),
		.in_data_21(config_reg_21_O),
		.in_data_22(ZextWrapper_20_32_inst1$self_O_in),
		.in_data_23(config_reg_23_O),
		.in_data_24(config_reg_24_O),
		.in_data_25(config_reg_25_O),
		.in_data_26(ZextWrapper_17_32_inst3$self_O_in),
		.in_data_27(config_reg_27_O),
		.in_data_28(config_reg_28_O),
		.in_data_29(config_reg_29_O),
		.in_data_3(ZextWrapper_17_32_inst0$self_O_in),
		.in_data_30(ZextWrapper_17_32_inst4$self_O_in),
		.in_data_31(config_reg_31_O),
		.in_data_32(config_reg_32_O),
		.in_data_33(config_reg_33_O),
		.in_data_34(ZextWrapper_20_32_inst2$self_O_in),
		.in_data_35(config_reg_35_O),
		.in_data_36(config_reg_36_O),
		.in_data_37(ZextWrapper_20_32_inst3$self_O_in),
		.in_data_38(config_reg_38_O),
		.in_data_39(config_reg_39_O),
		.in_data_4(config_reg_4_O),
		.in_data_40(config_reg_40_O),
		.in_data_41(ZextWrapper_25_32_inst0$self_O_in),
		.in_data_42(config_reg_42_O),
		.in_data_43(config_reg_43_O),
		.in_data_44(config_reg_44_O),
		.in_data_45(config_reg_45_O),
		.in_data_46(config_reg_46_O),
		.in_data_47(config_reg_47_O),
		.in_data_48(ZextWrapper_28_32_inst0$self_O_in),
		.in_data_49(config_reg_49_O),
		.in_data_5(config_reg_5_O),
		.in_data_50(config_reg_50_O),
		.in_data_51(ZextWrapper_20_32_inst4$self_O_in),
		.in_data_52(config_reg_52_O),
		.in_data_53(config_reg_53_O),
		.in_data_54(config_reg_54_O),
		.in_data_55(ZextWrapper_17_32_inst5$self_O_in),
		.in_data_56(config_reg_56_O),
		.in_data_57(config_reg_57_O),
		.in_data_58(config_reg_58_O),
		.in_data_59(ZextWrapper_17_32_inst6$self_O_in),
		.in_data_6(config_reg_6_O),
		.in_data_60(config_reg_60_O),
		.in_data_61(config_reg_61_O),
		.in_data_62(config_reg_62_O),
		.in_data_63(ZextWrapper_20_32_inst5$self_O_in),
		.in_data_64(config_reg_64_O),
		.in_data_65(config_reg_65_O),
		.in_data_66(ZextWrapper_20_32_inst6$self_O_in),
		.in_data_67(config_reg_67_O),
		.in_data_68(config_reg_68_O),
		.in_data_69(config_reg_69_O),
		.in_data_7(config_reg_7_O),
		.in_data_70(config_reg_70_O),
		.in_data_71(ZextWrapper_25_32_inst1$self_O_in),
		.in_data_72(config_reg_72_O),
		.in_data_73(config_reg_73_O),
		.in_data_74(config_reg_74_O),
		.in_data_75(ZextWrapper_17_32_inst7$self_O_in),
		.in_data_76(config_reg_76_O),
		.in_data_77(config_reg_77_O),
		.in_data_78(config_reg_78_O),
		.in_data_79(config_reg_79_O),
		.in_data_8(config_reg_8_O),
		.in_data_80(config_reg_80_O),
		.in_data_81(ZextWrapper_11_32_inst0$self_O_in),
		.in_data_9(config_reg_9_O),
		.in_sel(MuxWrapper_82_32_inst0_S_in),
		.out(MuxWrapper_82_32_inst0$Mux82xBits32_inst0$coreir_commonlib_mux82x32_inst0_out)
	);
	mantle_wire__typeBitIn7 MuxWrapper_82_32_inst0_S(
		.in(MuxWrapper_82_32_inst0_S_in),
		.out(self_config_config_addr_out[6:0])
	);
	coreir_or #(.width(1)) OR_CONFIG_EN_SRAM_0(
		.in0(config_1_write),
		.in1(config_1_read),
		.out(OR_CONFIG_EN_SRAM_0_out)
	);
	coreir_orr #(.width(1)) OR_CONFIG_RD_SRAM$orr_inst0(
		.in(config_1_write),
		.out(OR_CONFIG_RD_SRAM$orr_inst0_out)
	);
	coreir_orr #(.width(1)) OR_CONFIG_WR_SRAM$orr_inst0(
		.in(config_1_read),
		.out(OR_CONFIG_WR_SRAM$orr_inst0_out)
	);
	coreir_or #(.width(8)) OR_config_addr_FEATURE(
		.in0(config_config_addr),
		.in1(config_1_config_addr),
		.out(OR_config_addr_FEATURE_out)
	);
	coreir_or #(.width(32)) OR_config_data_FEATURE(
		.in0(config_config_data),
		.in1(config_1_config_data),
		.out(OR_config_data_FEATURE_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_11_32_inst0$bit_const_0_None(.out(ZextWrapper_11_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit11 ZextWrapper_11_32_inst0$self_I(
		.in(config_reg_81_O),
		.out(ZextWrapper_11_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_11_32_inst0$self_O_out;
	assign ZextWrapper_11_32_inst0$self_O_out = {ZextWrapper_11_32_inst0$bit_const_0_None_out, ZextWrapper_11_32_inst0$bit_const_0_None_out, ZextWrapper_11_32_inst0$bit_const_0_None_out, ZextWrapper_11_32_inst0$bit_const_0_None_out, ZextWrapper_11_32_inst0$bit_const_0_None_out, ZextWrapper_11_32_inst0$bit_const_0_None_out, ZextWrapper_11_32_inst0$bit_const_0_None_out, ZextWrapper_11_32_inst0$bit_const_0_None_out, ZextWrapper_11_32_inst0$bit_const_0_None_out, ZextWrapper_11_32_inst0$bit_const_0_None_out, ZextWrapper_11_32_inst0$bit_const_0_None_out, ZextWrapper_11_32_inst0$bit_const_0_None_out, ZextWrapper_11_32_inst0$bit_const_0_None_out, ZextWrapper_11_32_inst0$bit_const_0_None_out, ZextWrapper_11_32_inst0$bit_const_0_None_out, ZextWrapper_11_32_inst0$bit_const_0_None_out, ZextWrapper_11_32_inst0$bit_const_0_None_out, ZextWrapper_11_32_inst0$bit_const_0_None_out, ZextWrapper_11_32_inst0$bit_const_0_None_out, ZextWrapper_11_32_inst0$bit_const_0_None_out, ZextWrapper_11_32_inst0$bit_const_0_None_out, ZextWrapper_11_32_inst0$self_I_out[10:0]};
	mantle_wire__typeBitIn32 ZextWrapper_11_32_inst0$self_O(
		.in(ZextWrapper_11_32_inst0$self_O_in),
		.out(ZextWrapper_11_32_inst0$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_17_32_inst0$bit_const_0_None(.out(ZextWrapper_17_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit17 ZextWrapper_17_32_inst0$self_I(
		.in(config_reg_3_O),
		.out(ZextWrapper_17_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_17_32_inst0$self_O_out;
	assign ZextWrapper_17_32_inst0$self_O_out = {ZextWrapper_17_32_inst0$bit_const_0_None_out, ZextWrapper_17_32_inst0$bit_const_0_None_out, ZextWrapper_17_32_inst0$bit_const_0_None_out, ZextWrapper_17_32_inst0$bit_const_0_None_out, ZextWrapper_17_32_inst0$bit_const_0_None_out, ZextWrapper_17_32_inst0$bit_const_0_None_out, ZextWrapper_17_32_inst0$bit_const_0_None_out, ZextWrapper_17_32_inst0$bit_const_0_None_out, ZextWrapper_17_32_inst0$bit_const_0_None_out, ZextWrapper_17_32_inst0$bit_const_0_None_out, ZextWrapper_17_32_inst0$bit_const_0_None_out, ZextWrapper_17_32_inst0$bit_const_0_None_out, ZextWrapper_17_32_inst0$bit_const_0_None_out, ZextWrapper_17_32_inst0$bit_const_0_None_out, ZextWrapper_17_32_inst0$bit_const_0_None_out, ZextWrapper_17_32_inst0$self_I_out[16:0]};
	mantle_wire__typeBitIn32 ZextWrapper_17_32_inst0$self_O(
		.in(ZextWrapper_17_32_inst0$self_O_in),
		.out(ZextWrapper_17_32_inst0$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_17_32_inst1$bit_const_0_None(.out(ZextWrapper_17_32_inst1$bit_const_0_None_out));
	mantle_wire__typeBit17 ZextWrapper_17_32_inst1$self_I(
		.in(config_reg_11_O),
		.out(ZextWrapper_17_32_inst1$self_I_out)
	);
	wire [31:0] ZextWrapper_17_32_inst1$self_O_out;
	assign ZextWrapper_17_32_inst1$self_O_out = {ZextWrapper_17_32_inst1$bit_const_0_None_out, ZextWrapper_17_32_inst1$bit_const_0_None_out, ZextWrapper_17_32_inst1$bit_const_0_None_out, ZextWrapper_17_32_inst1$bit_const_0_None_out, ZextWrapper_17_32_inst1$bit_const_0_None_out, ZextWrapper_17_32_inst1$bit_const_0_None_out, ZextWrapper_17_32_inst1$bit_const_0_None_out, ZextWrapper_17_32_inst1$bit_const_0_None_out, ZextWrapper_17_32_inst1$bit_const_0_None_out, ZextWrapper_17_32_inst1$bit_const_0_None_out, ZextWrapper_17_32_inst1$bit_const_0_None_out, ZextWrapper_17_32_inst1$bit_const_0_None_out, ZextWrapper_17_32_inst1$bit_const_0_None_out, ZextWrapper_17_32_inst1$bit_const_0_None_out, ZextWrapper_17_32_inst1$bit_const_0_None_out, ZextWrapper_17_32_inst1$self_I_out[16:0]};
	mantle_wire__typeBitIn32 ZextWrapper_17_32_inst1$self_O(
		.in(ZextWrapper_17_32_inst1$self_O_in),
		.out(ZextWrapper_17_32_inst1$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_17_32_inst2$bit_const_0_None(.out(ZextWrapper_17_32_inst2$bit_const_0_None_out));
	mantle_wire__typeBit17 ZextWrapper_17_32_inst2$self_I(
		.in(config_reg_15_O),
		.out(ZextWrapper_17_32_inst2$self_I_out)
	);
	wire [31:0] ZextWrapper_17_32_inst2$self_O_out;
	assign ZextWrapper_17_32_inst2$self_O_out = {ZextWrapper_17_32_inst2$bit_const_0_None_out, ZextWrapper_17_32_inst2$bit_const_0_None_out, ZextWrapper_17_32_inst2$bit_const_0_None_out, ZextWrapper_17_32_inst2$bit_const_0_None_out, ZextWrapper_17_32_inst2$bit_const_0_None_out, ZextWrapper_17_32_inst2$bit_const_0_None_out, ZextWrapper_17_32_inst2$bit_const_0_None_out, ZextWrapper_17_32_inst2$bit_const_0_None_out, ZextWrapper_17_32_inst2$bit_const_0_None_out, ZextWrapper_17_32_inst2$bit_const_0_None_out, ZextWrapper_17_32_inst2$bit_const_0_None_out, ZextWrapper_17_32_inst2$bit_const_0_None_out, ZextWrapper_17_32_inst2$bit_const_0_None_out, ZextWrapper_17_32_inst2$bit_const_0_None_out, ZextWrapper_17_32_inst2$bit_const_0_None_out, ZextWrapper_17_32_inst2$self_I_out[16:0]};
	mantle_wire__typeBitIn32 ZextWrapper_17_32_inst2$self_O(
		.in(ZextWrapper_17_32_inst2$self_O_in),
		.out(ZextWrapper_17_32_inst2$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_17_32_inst3$bit_const_0_None(.out(ZextWrapper_17_32_inst3$bit_const_0_None_out));
	mantle_wire__typeBit17 ZextWrapper_17_32_inst3$self_I(
		.in(config_reg_26_O),
		.out(ZextWrapper_17_32_inst3$self_I_out)
	);
	wire [31:0] ZextWrapper_17_32_inst3$self_O_out;
	assign ZextWrapper_17_32_inst3$self_O_out = {ZextWrapper_17_32_inst3$bit_const_0_None_out, ZextWrapper_17_32_inst3$bit_const_0_None_out, ZextWrapper_17_32_inst3$bit_const_0_None_out, ZextWrapper_17_32_inst3$bit_const_0_None_out, ZextWrapper_17_32_inst3$bit_const_0_None_out, ZextWrapper_17_32_inst3$bit_const_0_None_out, ZextWrapper_17_32_inst3$bit_const_0_None_out, ZextWrapper_17_32_inst3$bit_const_0_None_out, ZextWrapper_17_32_inst3$bit_const_0_None_out, ZextWrapper_17_32_inst3$bit_const_0_None_out, ZextWrapper_17_32_inst3$bit_const_0_None_out, ZextWrapper_17_32_inst3$bit_const_0_None_out, ZextWrapper_17_32_inst3$bit_const_0_None_out, ZextWrapper_17_32_inst3$bit_const_0_None_out, ZextWrapper_17_32_inst3$bit_const_0_None_out, ZextWrapper_17_32_inst3$self_I_out[16:0]};
	mantle_wire__typeBitIn32 ZextWrapper_17_32_inst3$self_O(
		.in(ZextWrapper_17_32_inst3$self_O_in),
		.out(ZextWrapper_17_32_inst3$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_17_32_inst4$bit_const_0_None(.out(ZextWrapper_17_32_inst4$bit_const_0_None_out));
	mantle_wire__typeBit17 ZextWrapper_17_32_inst4$self_I(
		.in(config_reg_30_O),
		.out(ZextWrapper_17_32_inst4$self_I_out)
	);
	wire [31:0] ZextWrapper_17_32_inst4$self_O_out;
	assign ZextWrapper_17_32_inst4$self_O_out = {ZextWrapper_17_32_inst4$bit_const_0_None_out, ZextWrapper_17_32_inst4$bit_const_0_None_out, ZextWrapper_17_32_inst4$bit_const_0_None_out, ZextWrapper_17_32_inst4$bit_const_0_None_out, ZextWrapper_17_32_inst4$bit_const_0_None_out, ZextWrapper_17_32_inst4$bit_const_0_None_out, ZextWrapper_17_32_inst4$bit_const_0_None_out, ZextWrapper_17_32_inst4$bit_const_0_None_out, ZextWrapper_17_32_inst4$bit_const_0_None_out, ZextWrapper_17_32_inst4$bit_const_0_None_out, ZextWrapper_17_32_inst4$bit_const_0_None_out, ZextWrapper_17_32_inst4$bit_const_0_None_out, ZextWrapper_17_32_inst4$bit_const_0_None_out, ZextWrapper_17_32_inst4$bit_const_0_None_out, ZextWrapper_17_32_inst4$bit_const_0_None_out, ZextWrapper_17_32_inst4$self_I_out[16:0]};
	mantle_wire__typeBitIn32 ZextWrapper_17_32_inst4$self_O(
		.in(ZextWrapper_17_32_inst4$self_O_in),
		.out(ZextWrapper_17_32_inst4$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_17_32_inst5$bit_const_0_None(.out(ZextWrapper_17_32_inst5$bit_const_0_None_out));
	mantle_wire__typeBit17 ZextWrapper_17_32_inst5$self_I(
		.in(config_reg_55_O),
		.out(ZextWrapper_17_32_inst5$self_I_out)
	);
	wire [31:0] ZextWrapper_17_32_inst5$self_O_out;
	assign ZextWrapper_17_32_inst5$self_O_out = {ZextWrapper_17_32_inst5$bit_const_0_None_out, ZextWrapper_17_32_inst5$bit_const_0_None_out, ZextWrapper_17_32_inst5$bit_const_0_None_out, ZextWrapper_17_32_inst5$bit_const_0_None_out, ZextWrapper_17_32_inst5$bit_const_0_None_out, ZextWrapper_17_32_inst5$bit_const_0_None_out, ZextWrapper_17_32_inst5$bit_const_0_None_out, ZextWrapper_17_32_inst5$bit_const_0_None_out, ZextWrapper_17_32_inst5$bit_const_0_None_out, ZextWrapper_17_32_inst5$bit_const_0_None_out, ZextWrapper_17_32_inst5$bit_const_0_None_out, ZextWrapper_17_32_inst5$bit_const_0_None_out, ZextWrapper_17_32_inst5$bit_const_0_None_out, ZextWrapper_17_32_inst5$bit_const_0_None_out, ZextWrapper_17_32_inst5$bit_const_0_None_out, ZextWrapper_17_32_inst5$self_I_out[16:0]};
	mantle_wire__typeBitIn32 ZextWrapper_17_32_inst5$self_O(
		.in(ZextWrapper_17_32_inst5$self_O_in),
		.out(ZextWrapper_17_32_inst5$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_17_32_inst6$bit_const_0_None(.out(ZextWrapper_17_32_inst6$bit_const_0_None_out));
	mantle_wire__typeBit17 ZextWrapper_17_32_inst6$self_I(
		.in(config_reg_59_O),
		.out(ZextWrapper_17_32_inst6$self_I_out)
	);
	wire [31:0] ZextWrapper_17_32_inst6$self_O_out;
	assign ZextWrapper_17_32_inst6$self_O_out = {ZextWrapper_17_32_inst6$bit_const_0_None_out, ZextWrapper_17_32_inst6$bit_const_0_None_out, ZextWrapper_17_32_inst6$bit_const_0_None_out, ZextWrapper_17_32_inst6$bit_const_0_None_out, ZextWrapper_17_32_inst6$bit_const_0_None_out, ZextWrapper_17_32_inst6$bit_const_0_None_out, ZextWrapper_17_32_inst6$bit_const_0_None_out, ZextWrapper_17_32_inst6$bit_const_0_None_out, ZextWrapper_17_32_inst6$bit_const_0_None_out, ZextWrapper_17_32_inst6$bit_const_0_None_out, ZextWrapper_17_32_inst6$bit_const_0_None_out, ZextWrapper_17_32_inst6$bit_const_0_None_out, ZextWrapper_17_32_inst6$bit_const_0_None_out, ZextWrapper_17_32_inst6$bit_const_0_None_out, ZextWrapper_17_32_inst6$bit_const_0_None_out, ZextWrapper_17_32_inst6$self_I_out[16:0]};
	mantle_wire__typeBitIn32 ZextWrapper_17_32_inst6$self_O(
		.in(ZextWrapper_17_32_inst6$self_O_in),
		.out(ZextWrapper_17_32_inst6$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_17_32_inst7$bit_const_0_None(.out(ZextWrapper_17_32_inst7$bit_const_0_None_out));
	mantle_wire__typeBit17 ZextWrapper_17_32_inst7$self_I(
		.in(config_reg_75_O),
		.out(ZextWrapper_17_32_inst7$self_I_out)
	);
	wire [31:0] ZextWrapper_17_32_inst7$self_O_out;
	assign ZextWrapper_17_32_inst7$self_O_out = {ZextWrapper_17_32_inst7$bit_const_0_None_out, ZextWrapper_17_32_inst7$bit_const_0_None_out, ZextWrapper_17_32_inst7$bit_const_0_None_out, ZextWrapper_17_32_inst7$bit_const_0_None_out, ZextWrapper_17_32_inst7$bit_const_0_None_out, ZextWrapper_17_32_inst7$bit_const_0_None_out, ZextWrapper_17_32_inst7$bit_const_0_None_out, ZextWrapper_17_32_inst7$bit_const_0_None_out, ZextWrapper_17_32_inst7$bit_const_0_None_out, ZextWrapper_17_32_inst7$bit_const_0_None_out, ZextWrapper_17_32_inst7$bit_const_0_None_out, ZextWrapper_17_32_inst7$bit_const_0_None_out, ZextWrapper_17_32_inst7$bit_const_0_None_out, ZextWrapper_17_32_inst7$bit_const_0_None_out, ZextWrapper_17_32_inst7$bit_const_0_None_out, ZextWrapper_17_32_inst7$self_I_out[16:0]};
	mantle_wire__typeBitIn32 ZextWrapper_17_32_inst7$self_O(
		.in(ZextWrapper_17_32_inst7$self_O_in),
		.out(ZextWrapper_17_32_inst7$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_20_32_inst0$bit_const_0_None(.out(ZextWrapper_20_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit20 ZextWrapper_20_32_inst0$self_I(
		.in(config_reg_19_O),
		.out(ZextWrapper_20_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_20_32_inst0$self_O_out;
	assign ZextWrapper_20_32_inst0$self_O_out = {ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$bit_const_0_None_out, ZextWrapper_20_32_inst0$self_I_out[19:0]};
	mantle_wire__typeBitIn32 ZextWrapper_20_32_inst0$self_O(
		.in(ZextWrapper_20_32_inst0$self_O_in),
		.out(ZextWrapper_20_32_inst0$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_20_32_inst1$bit_const_0_None(.out(ZextWrapper_20_32_inst1$bit_const_0_None_out));
	mantle_wire__typeBit20 ZextWrapper_20_32_inst1$self_I(
		.in(config_reg_22_O),
		.out(ZextWrapper_20_32_inst1$self_I_out)
	);
	wire [31:0] ZextWrapper_20_32_inst1$self_O_out;
	assign ZextWrapper_20_32_inst1$self_O_out = {ZextWrapper_20_32_inst1$bit_const_0_None_out, ZextWrapper_20_32_inst1$bit_const_0_None_out, ZextWrapper_20_32_inst1$bit_const_0_None_out, ZextWrapper_20_32_inst1$bit_const_0_None_out, ZextWrapper_20_32_inst1$bit_const_0_None_out, ZextWrapper_20_32_inst1$bit_const_0_None_out, ZextWrapper_20_32_inst1$bit_const_0_None_out, ZextWrapper_20_32_inst1$bit_const_0_None_out, ZextWrapper_20_32_inst1$bit_const_0_None_out, ZextWrapper_20_32_inst1$bit_const_0_None_out, ZextWrapper_20_32_inst1$bit_const_0_None_out, ZextWrapper_20_32_inst1$bit_const_0_None_out, ZextWrapper_20_32_inst1$self_I_out[19:0]};
	mantle_wire__typeBitIn32 ZextWrapper_20_32_inst1$self_O(
		.in(ZextWrapper_20_32_inst1$self_O_in),
		.out(ZextWrapper_20_32_inst1$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_20_32_inst2$bit_const_0_None(.out(ZextWrapper_20_32_inst2$bit_const_0_None_out));
	mantle_wire__typeBit20 ZextWrapper_20_32_inst2$self_I(
		.in(config_reg_34_O),
		.out(ZextWrapper_20_32_inst2$self_I_out)
	);
	wire [31:0] ZextWrapper_20_32_inst2$self_O_out;
	assign ZextWrapper_20_32_inst2$self_O_out = {ZextWrapper_20_32_inst2$bit_const_0_None_out, ZextWrapper_20_32_inst2$bit_const_0_None_out, ZextWrapper_20_32_inst2$bit_const_0_None_out, ZextWrapper_20_32_inst2$bit_const_0_None_out, ZextWrapper_20_32_inst2$bit_const_0_None_out, ZextWrapper_20_32_inst2$bit_const_0_None_out, ZextWrapper_20_32_inst2$bit_const_0_None_out, ZextWrapper_20_32_inst2$bit_const_0_None_out, ZextWrapper_20_32_inst2$bit_const_0_None_out, ZextWrapper_20_32_inst2$bit_const_0_None_out, ZextWrapper_20_32_inst2$bit_const_0_None_out, ZextWrapper_20_32_inst2$bit_const_0_None_out, ZextWrapper_20_32_inst2$self_I_out[19:0]};
	mantle_wire__typeBitIn32 ZextWrapper_20_32_inst2$self_O(
		.in(ZextWrapper_20_32_inst2$self_O_in),
		.out(ZextWrapper_20_32_inst2$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_20_32_inst3$bit_const_0_None(.out(ZextWrapper_20_32_inst3$bit_const_0_None_out));
	mantle_wire__typeBit20 ZextWrapper_20_32_inst3$self_I(
		.in(config_reg_37_O),
		.out(ZextWrapper_20_32_inst3$self_I_out)
	);
	wire [31:0] ZextWrapper_20_32_inst3$self_O_out;
	assign ZextWrapper_20_32_inst3$self_O_out = {ZextWrapper_20_32_inst3$bit_const_0_None_out, ZextWrapper_20_32_inst3$bit_const_0_None_out, ZextWrapper_20_32_inst3$bit_const_0_None_out, ZextWrapper_20_32_inst3$bit_const_0_None_out, ZextWrapper_20_32_inst3$bit_const_0_None_out, ZextWrapper_20_32_inst3$bit_const_0_None_out, ZextWrapper_20_32_inst3$bit_const_0_None_out, ZextWrapper_20_32_inst3$bit_const_0_None_out, ZextWrapper_20_32_inst3$bit_const_0_None_out, ZextWrapper_20_32_inst3$bit_const_0_None_out, ZextWrapper_20_32_inst3$bit_const_0_None_out, ZextWrapper_20_32_inst3$bit_const_0_None_out, ZextWrapper_20_32_inst3$self_I_out[19:0]};
	mantle_wire__typeBitIn32 ZextWrapper_20_32_inst3$self_O(
		.in(ZextWrapper_20_32_inst3$self_O_in),
		.out(ZextWrapper_20_32_inst3$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_20_32_inst4$bit_const_0_None(.out(ZextWrapper_20_32_inst4$bit_const_0_None_out));
	mantle_wire__typeBit20 ZextWrapper_20_32_inst4$self_I(
		.in(config_reg_51_O),
		.out(ZextWrapper_20_32_inst4$self_I_out)
	);
	wire [31:0] ZextWrapper_20_32_inst4$self_O_out;
	assign ZextWrapper_20_32_inst4$self_O_out = {ZextWrapper_20_32_inst4$bit_const_0_None_out, ZextWrapper_20_32_inst4$bit_const_0_None_out, ZextWrapper_20_32_inst4$bit_const_0_None_out, ZextWrapper_20_32_inst4$bit_const_0_None_out, ZextWrapper_20_32_inst4$bit_const_0_None_out, ZextWrapper_20_32_inst4$bit_const_0_None_out, ZextWrapper_20_32_inst4$bit_const_0_None_out, ZextWrapper_20_32_inst4$bit_const_0_None_out, ZextWrapper_20_32_inst4$bit_const_0_None_out, ZextWrapper_20_32_inst4$bit_const_0_None_out, ZextWrapper_20_32_inst4$bit_const_0_None_out, ZextWrapper_20_32_inst4$bit_const_0_None_out, ZextWrapper_20_32_inst4$self_I_out[19:0]};
	mantle_wire__typeBitIn32 ZextWrapper_20_32_inst4$self_O(
		.in(ZextWrapper_20_32_inst4$self_O_in),
		.out(ZextWrapper_20_32_inst4$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_20_32_inst5$bit_const_0_None(.out(ZextWrapper_20_32_inst5$bit_const_0_None_out));
	mantle_wire__typeBit20 ZextWrapper_20_32_inst5$self_I(
		.in(config_reg_63_O),
		.out(ZextWrapper_20_32_inst5$self_I_out)
	);
	wire [31:0] ZextWrapper_20_32_inst5$self_O_out;
	assign ZextWrapper_20_32_inst5$self_O_out = {ZextWrapper_20_32_inst5$bit_const_0_None_out, ZextWrapper_20_32_inst5$bit_const_0_None_out, ZextWrapper_20_32_inst5$bit_const_0_None_out, ZextWrapper_20_32_inst5$bit_const_0_None_out, ZextWrapper_20_32_inst5$bit_const_0_None_out, ZextWrapper_20_32_inst5$bit_const_0_None_out, ZextWrapper_20_32_inst5$bit_const_0_None_out, ZextWrapper_20_32_inst5$bit_const_0_None_out, ZextWrapper_20_32_inst5$bit_const_0_None_out, ZextWrapper_20_32_inst5$bit_const_0_None_out, ZextWrapper_20_32_inst5$bit_const_0_None_out, ZextWrapper_20_32_inst5$bit_const_0_None_out, ZextWrapper_20_32_inst5$self_I_out[19:0]};
	mantle_wire__typeBitIn32 ZextWrapper_20_32_inst5$self_O(
		.in(ZextWrapper_20_32_inst5$self_O_in),
		.out(ZextWrapper_20_32_inst5$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_20_32_inst6$bit_const_0_None(.out(ZextWrapper_20_32_inst6$bit_const_0_None_out));
	mantle_wire__typeBit20 ZextWrapper_20_32_inst6$self_I(
		.in(config_reg_66_O),
		.out(ZextWrapper_20_32_inst6$self_I_out)
	);
	wire [31:0] ZextWrapper_20_32_inst6$self_O_out;
	assign ZextWrapper_20_32_inst6$self_O_out = {ZextWrapper_20_32_inst6$bit_const_0_None_out, ZextWrapper_20_32_inst6$bit_const_0_None_out, ZextWrapper_20_32_inst6$bit_const_0_None_out, ZextWrapper_20_32_inst6$bit_const_0_None_out, ZextWrapper_20_32_inst6$bit_const_0_None_out, ZextWrapper_20_32_inst6$bit_const_0_None_out, ZextWrapper_20_32_inst6$bit_const_0_None_out, ZextWrapper_20_32_inst6$bit_const_0_None_out, ZextWrapper_20_32_inst6$bit_const_0_None_out, ZextWrapper_20_32_inst6$bit_const_0_None_out, ZextWrapper_20_32_inst6$bit_const_0_None_out, ZextWrapper_20_32_inst6$bit_const_0_None_out, ZextWrapper_20_32_inst6$self_I_out[19:0]};
	mantle_wire__typeBitIn32 ZextWrapper_20_32_inst6$self_O(
		.in(ZextWrapper_20_32_inst6$self_O_in),
		.out(ZextWrapper_20_32_inst6$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_25_32_inst0$bit_const_0_None(.out(ZextWrapper_25_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit25 ZextWrapper_25_32_inst0$self_I(
		.in(config_reg_41_O),
		.out(ZextWrapper_25_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_25_32_inst0$self_O_out;
	assign ZextWrapper_25_32_inst0$self_O_out = {ZextWrapper_25_32_inst0$bit_const_0_None_out, ZextWrapper_25_32_inst0$bit_const_0_None_out, ZextWrapper_25_32_inst0$bit_const_0_None_out, ZextWrapper_25_32_inst0$bit_const_0_None_out, ZextWrapper_25_32_inst0$bit_const_0_None_out, ZextWrapper_25_32_inst0$bit_const_0_None_out, ZextWrapper_25_32_inst0$bit_const_0_None_out, ZextWrapper_25_32_inst0$self_I_out[24:0]};
	mantle_wire__typeBitIn32 ZextWrapper_25_32_inst0$self_O(
		.in(ZextWrapper_25_32_inst0$self_O_in),
		.out(ZextWrapper_25_32_inst0$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_25_32_inst1$bit_const_0_None(.out(ZextWrapper_25_32_inst1$bit_const_0_None_out));
	mantle_wire__typeBit25 ZextWrapper_25_32_inst1$self_I(
		.in(config_reg_71_O),
		.out(ZextWrapper_25_32_inst1$self_I_out)
	);
	wire [31:0] ZextWrapper_25_32_inst1$self_O_out;
	assign ZextWrapper_25_32_inst1$self_O_out = {ZextWrapper_25_32_inst1$bit_const_0_None_out, ZextWrapper_25_32_inst1$bit_const_0_None_out, ZextWrapper_25_32_inst1$bit_const_0_None_out, ZextWrapper_25_32_inst1$bit_const_0_None_out, ZextWrapper_25_32_inst1$bit_const_0_None_out, ZextWrapper_25_32_inst1$bit_const_0_None_out, ZextWrapper_25_32_inst1$bit_const_0_None_out, ZextWrapper_25_32_inst1$self_I_out[24:0]};
	mantle_wire__typeBitIn32 ZextWrapper_25_32_inst1$self_O(
		.in(ZextWrapper_25_32_inst1$self_O_in),
		.out(ZextWrapper_25_32_inst1$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_26_32_inst0$bit_const_0_None(.out(ZextWrapper_26_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit26 ZextWrapper_26_32_inst0$self_I(
		.in(config_reg_0_O),
		.out(ZextWrapper_26_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_26_32_inst0$self_O_out;
	assign ZextWrapper_26_32_inst0$self_O_out = {ZextWrapper_26_32_inst0$bit_const_0_None_out, ZextWrapper_26_32_inst0$bit_const_0_None_out, ZextWrapper_26_32_inst0$bit_const_0_None_out, ZextWrapper_26_32_inst0$bit_const_0_None_out, ZextWrapper_26_32_inst0$bit_const_0_None_out, ZextWrapper_26_32_inst0$bit_const_0_None_out, ZextWrapper_26_32_inst0$self_I_out[25:0]};
	mantle_wire__typeBitIn32 ZextWrapper_26_32_inst0$self_O(
		.in(ZextWrapper_26_32_inst0$self_O_in),
		.out(ZextWrapper_26_32_inst0$self_O_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_28_32_inst0$bit_const_0_None(.out(ZextWrapper_28_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit28 ZextWrapper_28_32_inst0$self_I(
		.in(config_reg_48_O),
		.out(ZextWrapper_28_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_28_32_inst0$self_O_out;
	assign ZextWrapper_28_32_inst0$self_O_out = {ZextWrapper_28_32_inst0$bit_const_0_None_out, ZextWrapper_28_32_inst0$bit_const_0_None_out, ZextWrapper_28_32_inst0$bit_const_0_None_out, ZextWrapper_28_32_inst0$bit_const_0_None_out, ZextWrapper_28_32_inst0$self_I_out[27:0]};
	mantle_wire__typeBitIn32 ZextWrapper_28_32_inst0$self_O(
		.in(ZextWrapper_28_32_inst0$self_O_in),
		.out(ZextWrapper_28_32_inst0$self_O_out)
	);
	ConfigRegister_26_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_1 config_reg_1(
		.clk(clk),
		.reset(reset),
		.O(config_reg_1_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_10 config_reg_10(
		.clk(clk),
		.reset(reset),
		.O(config_reg_10_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_17_8_32_11 config_reg_11(
		.clk(clk),
		.reset(reset),
		.O(config_reg_11_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_12 config_reg_12(
		.clk(clk),
		.reset(reset),
		.O(config_reg_12_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_13 config_reg_13(
		.clk(clk),
		.reset(reset),
		.O(config_reg_13_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_14 config_reg_14(
		.clk(clk),
		.reset(reset),
		.O(config_reg_14_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_17_8_32_15 config_reg_15(
		.clk(clk),
		.reset(reset),
		.O(config_reg_15_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_16 config_reg_16(
		.clk(clk),
		.reset(reset),
		.O(config_reg_16_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_17 config_reg_17(
		.clk(clk),
		.reset(reset),
		.O(config_reg_17_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_18 config_reg_18(
		.clk(clk),
		.reset(reset),
		.O(config_reg_18_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_20_8_32_19 config_reg_19(
		.clk(clk),
		.reset(reset),
		.O(config_reg_19_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_2 config_reg_2(
		.clk(clk),
		.reset(reset),
		.O(config_reg_2_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_20 config_reg_20(
		.clk(clk),
		.reset(reset),
		.O(config_reg_20_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_21 config_reg_21(
		.clk(clk),
		.reset(reset),
		.O(config_reg_21_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_20_8_32_22 config_reg_22(
		.clk(clk),
		.reset(reset),
		.O(config_reg_22_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_23 config_reg_23(
		.clk(clk),
		.reset(reset),
		.O(config_reg_23_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_24 config_reg_24(
		.clk(clk),
		.reset(reset),
		.O(config_reg_24_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_25 config_reg_25(
		.clk(clk),
		.reset(reset),
		.O(config_reg_25_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_17_8_32_26 config_reg_26(
		.clk(clk),
		.reset(reset),
		.O(config_reg_26_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_27 config_reg_27(
		.clk(clk),
		.reset(reset),
		.O(config_reg_27_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_28 config_reg_28(
		.clk(clk),
		.reset(reset),
		.O(config_reg_28_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_29 config_reg_29(
		.clk(clk),
		.reset(reset),
		.O(config_reg_29_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_17_8_32_3 config_reg_3(
		.clk(clk),
		.reset(reset),
		.O(config_reg_3_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_17_8_32_30 config_reg_30(
		.clk(clk),
		.reset(reset),
		.O(config_reg_30_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_31 config_reg_31(
		.clk(clk),
		.reset(reset),
		.O(config_reg_31_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_32 config_reg_32(
		.clk(clk),
		.reset(reset),
		.O(config_reg_32_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_33 config_reg_33(
		.clk(clk),
		.reset(reset),
		.O(config_reg_33_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_20_8_32_34 config_reg_34(
		.clk(clk),
		.reset(reset),
		.O(config_reg_34_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_35 config_reg_35(
		.clk(clk),
		.reset(reset),
		.O(config_reg_35_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_36 config_reg_36(
		.clk(clk),
		.reset(reset),
		.O(config_reg_36_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_20_8_32_37 config_reg_37(
		.clk(clk),
		.reset(reset),
		.O(config_reg_37_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_38 config_reg_38(
		.clk(clk),
		.reset(reset),
		.O(config_reg_38_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_39 config_reg_39(
		.clk(clk),
		.reset(reset),
		.O(config_reg_39_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_4 config_reg_4(
		.clk(clk),
		.reset(reset),
		.O(config_reg_4_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_40 config_reg_40(
		.clk(clk),
		.reset(reset),
		.O(config_reg_40_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_25_8_32_41 config_reg_41(
		.clk(clk),
		.reset(reset),
		.O(config_reg_41_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_42 config_reg_42(
		.clk(clk),
		.reset(reset),
		.O(config_reg_42_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_43 config_reg_43(
		.clk(clk),
		.reset(reset),
		.O(config_reg_43_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_44 config_reg_44(
		.clk(clk),
		.reset(reset),
		.O(config_reg_44_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_45 config_reg_45(
		.clk(clk),
		.reset(reset),
		.O(config_reg_45_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_46 config_reg_46(
		.clk(clk),
		.reset(reset),
		.O(config_reg_46_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_47 config_reg_47(
		.clk(clk),
		.reset(reset),
		.O(config_reg_47_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_28_8_32_48 config_reg_48(
		.clk(clk),
		.reset(reset),
		.O(config_reg_48_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_49 config_reg_49(
		.clk(clk),
		.reset(reset),
		.O(config_reg_49_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_5 config_reg_5(
		.clk(clk),
		.reset(reset),
		.O(config_reg_5_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_50 config_reg_50(
		.clk(clk),
		.reset(reset),
		.O(config_reg_50_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_20_8_32_51 config_reg_51(
		.clk(clk),
		.reset(reset),
		.O(config_reg_51_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_52 config_reg_52(
		.clk(clk),
		.reset(reset),
		.O(config_reg_52_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_53 config_reg_53(
		.clk(clk),
		.reset(reset),
		.O(config_reg_53_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_54 config_reg_54(
		.clk(clk),
		.reset(reset),
		.O(config_reg_54_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_17_8_32_55 config_reg_55(
		.clk(clk),
		.reset(reset),
		.O(config_reg_55_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_56 config_reg_56(
		.clk(clk),
		.reset(reset),
		.O(config_reg_56_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_57 config_reg_57(
		.clk(clk),
		.reset(reset),
		.O(config_reg_57_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_58 config_reg_58(
		.clk(clk),
		.reset(reset),
		.O(config_reg_58_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_17_8_32_59 config_reg_59(
		.clk(clk),
		.reset(reset),
		.O(config_reg_59_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_6 config_reg_6(
		.clk(clk),
		.reset(reset),
		.O(config_reg_6_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_60 config_reg_60(
		.clk(clk),
		.reset(reset),
		.O(config_reg_60_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_61 config_reg_61(
		.clk(clk),
		.reset(reset),
		.O(config_reg_61_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_62 config_reg_62(
		.clk(clk),
		.reset(reset),
		.O(config_reg_62_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_20_8_32_63 config_reg_63(
		.clk(clk),
		.reset(reset),
		.O(config_reg_63_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_64 config_reg_64(
		.clk(clk),
		.reset(reset),
		.O(config_reg_64_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_65 config_reg_65(
		.clk(clk),
		.reset(reset),
		.O(config_reg_65_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_20_8_32_66 config_reg_66(
		.clk(clk),
		.reset(reset),
		.O(config_reg_66_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_67 config_reg_67(
		.clk(clk),
		.reset(reset),
		.O(config_reg_67_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_68 config_reg_68(
		.clk(clk),
		.reset(reset),
		.O(config_reg_68_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_69 config_reg_69(
		.clk(clk),
		.reset(reset),
		.O(config_reg_69_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_7 config_reg_7(
		.clk(clk),
		.reset(reset),
		.O(config_reg_7_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_70 config_reg_70(
		.clk(clk),
		.reset(reset),
		.O(config_reg_70_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_25_8_32_71 config_reg_71(
		.clk(clk),
		.reset(reset),
		.O(config_reg_71_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_72 config_reg_72(
		.clk(clk),
		.reset(reset),
		.O(config_reg_72_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_73 config_reg_73(
		.clk(clk),
		.reset(reset),
		.O(config_reg_73_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_74 config_reg_74(
		.clk(clk),
		.reset(reset),
		.O(config_reg_74_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_17_8_32_75 config_reg_75(
		.clk(clk),
		.reset(reset),
		.O(config_reg_75_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_76 config_reg_76(
		.clk(clk),
		.reset(reset),
		.O(config_reg_76_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_77 config_reg_77(
		.clk(clk),
		.reset(reset),
		.O(config_reg_77_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_78 config_reg_78(
		.clk(clk),
		.reset(reset),
		.O(config_reg_78_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_79 config_reg_79(
		.clk(clk),
		.reset(reset),
		.O(config_reg_79_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_8 config_reg_8(
		.clk(clk),
		.reset(reset),
		.O(config_reg_8_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_80 config_reg_80(
		.clk(clk),
		.reset(reset),
		.O(config_reg_80_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_11_8_32_81 config_reg_81(
		.clk(clk),
		.reset(reset),
		.O(config_reg_81_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_9 config_reg_9(
		.clk(clk),
		.reset(reset),
		.O(config_reg_9_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	coreir_wrap coreir_wrapInAsyncReset_inst0(
		.in(reset),
		.out(coreir_wrapInAsyncReset_inst0_out)
	);
	coreir_wrap coreir_wrapOutAsyncReset_inst0(
		.in(Invert1_inst0_out[0]),
		.out(coreir_wrapOutAsyncReset_inst0_out)
	);
	flush_reg_sel flush_reg_sel_inst0(
		.I(config_reg_0_O),
		.O(flush_reg_sel_inst0_O)
	);
	flush_reg_value flush_reg_value_inst0(
		.I(config_reg_0_O),
		.O(flush_reg_value_inst0_O)
	);
	coreir_mux #(.width(1)) flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(flush),
		.in1(flush_reg_value_inst0_O),
		.sel(flush_reg_sel_inst0_O[0]),
		.out(flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	input_width_1_num_0_reg_sel input_width_1_num_0_reg_sel_inst0(
		.I(config_reg_0_O),
		.O(input_width_1_num_0_reg_sel_inst0_O)
	);
	input_width_1_num_0_reg_value input_width_1_num_0_reg_value_inst0(
		.I(config_reg_0_O),
		.O(input_width_1_num_0_reg_value_inst0_O)
	);
	coreir_mux #(.width(1)) input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(input_width_1_num_0),
		.in1(input_width_1_num_0_reg_value_inst0_O),
		.sel(input_width_1_num_0_reg_sel_inst0_O[0]),
		.out(input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	input_width_1_num_1_reg_sel input_width_1_num_1_reg_sel_inst0(
		.I(config_reg_0_O),
		.O(input_width_1_num_1_reg_sel_inst0_O)
	);
	input_width_1_num_1_reg_value input_width_1_num_1_reg_value_inst0(
		.I(config_reg_0_O),
		.O(input_width_1_num_1_reg_value_inst0_O)
	);
	coreir_mux #(.width(1)) input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(input_width_1_num_1),
		.in1(input_width_1_num_1_reg_value_inst0_O),
		.sel(input_width_1_num_1_reg_sel_inst0_O[0]),
		.out(input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality_inst0(
		.I(config_reg_0_O),
		.O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality_inst0_O)
	);
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0 mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0_inst0(
		.I(config_reg_0_O),
		.O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0_inst0_O)
	);
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1 mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1_inst0(
		.I(config_reg_1_O),
		.O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1_inst0_O)
	);
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2 mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2_inst0(
		.I(config_reg_1_O),
		.O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2_inst0_O)
	);
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3 mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3_inst0(
		.I(config_reg_2_O),
		.O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3_inst0_O)
	);
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4 mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4_inst0(
		.I(config_reg_2_O),
		.O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4_inst0_O)
	);
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5 mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5_inst0(
		.I(config_reg_3_O),
		.O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5_inst0_O)
	);
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable_inst0(
		.I(config_reg_3_O),
		.O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable_inst0_O)
	);
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr_inst0(
		.I(config_reg_4_O),
		.O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr_inst0_O)
	);
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0 mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0_inst0(
		.I(config_reg_4_O),
		.O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0_inst0_O)
	);
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1 mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1_inst0(
		.I(config_reg_5_O),
		.O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1_inst0_O)
	);
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2 mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2_inst0(
		.I(config_reg_5_O),
		.O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2_inst0_O)
	);
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3 mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3_inst0(
		.I(config_reg_6_O),
		.O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3_inst0_O)
	);
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4 mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4_inst0(
		.I(config_reg_6_O),
		.O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4_inst0_O)
	);
	mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5 mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5_inst0(
		.I(config_reg_7_O),
		.O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr_inst0(
		.I(config_reg_7_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_0_inst0(
		.I(config_reg_7_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_0_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_1_inst0(
		.I(config_reg_7_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_1_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_2_inst0(
		.I(config_reg_7_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_2_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_3_inst0(
		.I(config_reg_8_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_3_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_4_inst0(
		.I(config_reg_8_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_4_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_5_inst0(
		.I(config_reg_8_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_5_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr_inst0(
		.I(config_reg_8_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_0_inst0(
		.I(config_reg_8_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_0_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_1_inst0(
		.I(config_reg_8_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_1_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_2_inst0(
		.I(config_reg_8_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_2_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_3_inst0(
		.I(config_reg_8_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_3_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_4_inst0(
		.I(config_reg_9_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_4_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_5_inst0(
		.I(config_reg_9_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_5_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr_inst0(
		.I(config_reg_9_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0_inst0(
		.I(config_reg_9_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1_inst0(
		.I(config_reg_9_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2_inst0(
		.I(config_reg_9_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_3_inst0(
		.I(config_reg_9_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_3_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_4_inst0(
		.I(config_reg_9_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_4_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_5_inst0(
		.I(config_reg_10_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_5_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr_inst0(
		.I(config_reg_10_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0_inst0(
		.I(config_reg_10_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1_inst0(
		.I(config_reg_10_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2_inst0(
		.I(config_reg_10_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_3_inst0(
		.I(config_reg_10_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_3_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_4_inst0(
		.I(config_reg_10_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_4_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_5_inst0(
		.I(config_reg_10_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_5_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable_inst0(
		.I(config_reg_11_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr_inst0(
		.I(config_reg_11_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0_inst0(
		.I(config_reg_12_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1_inst0(
		.I(config_reg_12_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2_inst0(
		.I(config_reg_13_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3_inst0(
		.I(config_reg_13_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4_inst0(
		.I(config_reg_14_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5_inst0(
		.I(config_reg_14_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable_inst0(
		.I(config_reg_15_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr_inst0(
		.I(config_reg_15_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0_inst0(
		.I(config_reg_16_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1_inst0(
		.I(config_reg_16_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2_inst0(
		.I(config_reg_17_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3_inst0(
		.I(config_reg_17_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4_inst0(
		.I(config_reg_18_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5_inst0(
		.I(config_reg_18_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality_inst0(
		.I(config_reg_19_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0_inst0(
		.I(config_reg_19_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1_inst0(
		.I(config_reg_20_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2_inst0(
		.I(config_reg_20_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_3_inst0(
		.I(config_reg_21_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_3_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_4_inst0(
		.I(config_reg_21_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_4_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_5_inst0(
		.I(config_reg_22_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_5_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality_inst0(
		.I(config_reg_22_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0_inst0(
		.I(config_reg_23_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1_inst0(
		.I(config_reg_23_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2_inst0(
		.I(config_reg_24_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_3_inst0(
		.I(config_reg_24_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_3_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_4_inst0(
		.I(config_reg_25_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_4_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_5_inst0(
		.I(config_reg_25_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_5_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable_inst0(
		.I(config_reg_26_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr_inst0(
		.I(config_reg_26_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0_inst0(
		.I(config_reg_27_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1_inst0(
		.I(config_reg_27_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2_inst0(
		.I(config_reg_28_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3_inst0(
		.I(config_reg_28_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4_inst0(
		.I(config_reg_29_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5_inst0(
		.I(config_reg_29_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable_inst0(
		.I(config_reg_30_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr_inst0(
		.I(config_reg_30_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0_inst0(
		.I(config_reg_31_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1_inst0(
		.I(config_reg_31_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2_inst0(
		.I(config_reg_32_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3_inst0(
		.I(config_reg_32_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4_inst0(
		.I(config_reg_33_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5_inst0(
		.I(config_reg_33_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality_inst0(
		.I(config_reg_34_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0_inst0(
		.I(config_reg_34_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1_inst0(
		.I(config_reg_35_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2_inst0(
		.I(config_reg_35_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3_inst0(
		.I(config_reg_36_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4_inst0(
		.I(config_reg_36_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5_inst0(
		.I(config_reg_37_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality_inst0(
		.I(config_reg_37_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0_inst0(
		.I(config_reg_38_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1_inst0(
		.I(config_reg_38_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2_inst0(
		.I(config_reg_39_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3_inst0(
		.I(config_reg_39_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4_inst0(
		.I(config_reg_40_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5_inst0(
		.I(config_reg_40_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en_inst0(
		.I(config_reg_41_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr_inst0(
		.I(config_reg_41_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_0_inst0(
		.I(config_reg_41_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_0_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_1_inst0(
		.I(config_reg_41_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_1_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_2_inst0(
		.I(config_reg_42_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_2_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_3_inst0(
		.I(config_reg_42_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_3_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_4_inst0(
		.I(config_reg_42_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_4_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_5_inst0(
		.I(config_reg_42_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_5_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr_inst0(
		.I(config_reg_43_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_0_inst0(
		.I(config_reg_43_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_0_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_1_inst0(
		.I(config_reg_43_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_1_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_2_inst0(
		.I(config_reg_43_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_2_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_3_inst0(
		.I(config_reg_44_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_3_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_4_inst0(
		.I(config_reg_44_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_4_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_5_inst0(
		.I(config_reg_44_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_5_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr_inst0(
		.I(config_reg_44_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0_inst0(
		.I(config_reg_45_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1_inst0(
		.I(config_reg_45_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2_inst0(
		.I(config_reg_45_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3_inst0(
		.I(config_reg_45_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4_inst0(
		.I(config_reg_46_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5_inst0(
		.I(config_reg_46_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr_inst0(
		.I(config_reg_46_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0_inst0(
		.I(config_reg_46_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1_inst0(
		.I(config_reg_47_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2_inst0(
		.I(config_reg_47_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3_inst0(
		.I(config_reg_47_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4_inst0(
		.I(config_reg_47_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4_inst0_O)
	);
	mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5_inst0(
		.I(config_reg_48_O),
		.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5_inst0_O)
	);
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality_inst0(
	// 	.I(config_reg_48_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0_inst0(
	// 	.I(config_reg_48_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1_inst0(
	// 	.I(config_reg_49_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2_inst0(
	// 	.I(config_reg_49_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3_inst0(
	// 	.I(config_reg_50_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4_inst0(
	// 	.I(config_reg_50_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5_inst0(
	// 	.I(config_reg_51_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality_inst0(
	// 	.I(config_reg_51_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0_inst0(
	// 	.I(config_reg_52_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1_inst0(
	// 	.I(config_reg_52_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2_inst0(
	// 	.I(config_reg_53_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3_inst0(
	// 	.I(config_reg_53_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4_inst0(
	// 	.I(config_reg_54_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5_inst0(
	// 	.I(config_reg_54_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable_inst0(
	// 	.I(config_reg_55_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr_inst0(
	// 	.I(config_reg_55_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0_inst0(
	// 	.I(config_reg_56_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1_inst0(
	// 	.I(config_reg_56_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2_inst0(
	// 	.I(config_reg_57_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3_inst0(
	// 	.I(config_reg_57_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4_inst0(
	// 	.I(config_reg_58_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5_inst0(
	// 	.I(config_reg_58_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable_inst0(
	// 	.I(config_reg_59_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr_inst0(
	// 	.I(config_reg_59_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0_inst0(
	// 	.I(config_reg_60_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1_inst0(
	// 	.I(config_reg_60_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2_inst0(
	// 	.I(config_reg_61_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3_inst0(
	// 	.I(config_reg_61_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4_inst0(
	// 	.I(config_reg_62_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5_inst0(
	// 	.I(config_reg_62_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality_inst0(
	// 	.I(config_reg_63_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0_inst0(
	// 	.I(config_reg_63_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1_inst0(
	// 	.I(config_reg_64_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2_inst0(
	// 	.I(config_reg_64_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3_inst0(
	// 	.I(config_reg_65_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4_inst0(
	// 	.I(config_reg_65_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5_inst0(
	// 	.I(config_reg_66_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality_inst0(
	// 	.I(config_reg_66_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0_inst0(
	// 	.I(config_reg_67_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1_inst0(
	// 	.I(config_reg_67_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2_inst0(
	// 	.I(config_reg_68_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3_inst0(
	// 	.I(config_reg_68_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4_inst0(
	// 	.I(config_reg_69_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5_inst0(
	// 	.I(config_reg_69_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr_inst0(
	// 	.I(config_reg_70_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0_inst0(
	// 	.I(config_reg_70_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1_inst0(
	// 	.I(config_reg_70_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2_inst0(
	// 	.I(config_reg_70_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3_inst0(
	// 	.I(config_reg_70_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4_inst0(
	// 	.I(config_reg_70_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5_inst0(
	// 	.I(config_reg_70_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr_inst0(
	// 	.I(config_reg_70_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0_inst0(
	// 	.I(config_reg_71_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1_inst0(
	// 	.I(config_reg_71_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2_inst0(
	// 	.I(config_reg_71_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3_inst0(
	// 	.I(config_reg_71_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4_inst0(
	// 	.I(config_reg_71_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5_inst0(
	// 	.I(config_reg_71_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable_inst0(
	// 	.I(config_reg_71_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr_inst0(
	// 	.I(config_reg_72_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0_inst0(
	// 	.I(config_reg_72_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1_inst0(
	// 	.I(config_reg_73_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2_inst0(
	// 	.I(config_reg_73_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3_inst0(
	// 	.I(config_reg_74_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4_inst0(
	// 	.I(config_reg_74_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5_inst0(
	// 	.I(config_reg_75_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable_inst0(
	// 	.I(config_reg_75_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr_inst0(
	// 	.I(config_reg_76_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0_inst0(
	// 	.I(config_reg_76_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1_inst0(
	// 	.I(config_reg_77_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2_inst0(
	// 	.I(config_reg_77_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3_inst0(
	// 	.I(config_reg_78_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4_inst0(
	// 	.I(config_reg_78_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5_inst0(
	// 	.I(config_reg_79_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr_inst0(
	// 	.I(config_reg_79_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0_inst0(
	// 	.I(config_reg_79_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1_inst0(
	// 	.I(config_reg_79_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2_inst0(
	// 	.I(config_reg_79_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3_inst0(
	// 	.I(config_reg_80_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4_inst0(
	// 	.I(config_reg_80_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5_inst0(
	// 	.I(config_reg_80_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr_inst0(
	// 	.I(config_reg_80_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0_inst0(
	// 	.I(config_reg_80_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1_inst0(
	// 	.I(config_reg_80_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2_inst0(
	// 	.I(config_reg_80_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3_inst0(
	// 	.I(config_reg_80_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4_inst0(
	// 	.I(config_reg_81_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4_inst0_O)
	// );
	// mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5_inst0(
	// 	.I(config_reg_81_O),
	// 	.O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5_inst0_O)
	// );
	mode mode_inst0(
		.I(config_reg_81_O),
		.O(mode_inst0_O)
	);
	mantle_wire__typeBit8 self_config_config_addr(
		.in(config_config_addr),
		.out(self_config_config_addr_out)
	);
	tile_en tile_en_inst0(
		.I(config_reg_81_O),
		.O(tile_en_inst0_O)
	);
	assign output_width_16_num_0 = LakeTop_W_inst0_output_width_16_num_0;
	assign output_width_16_num_1 = LakeTop_W_inst0_output_width_16_num_1;
	assign output_width_1_num_0 = LakeTop_W_inst0_output_width_1_num_0;
	assign output_width_1_num_1 = LakeTop_W_inst0_output_width_1_num_1;
	assign output_width_1_num_2 = LakeTop_W_inst0_output_width_1_num_2;
	assign read_config_data = MuxWrapper_82_32_inst0$Mux82xBits32_inst0$coreir_commonlib_mux82x32_inst0_out;
	assign read_config_data_1 = LakeTop_W_inst0_config_data_out;
endmodule
module Cond (
	code,
	alu,
	lut,
	Z,
	N,
	C,
	V,
	O,
	CLK,
	ASYNCRESET
);
	input [4:0] code;
	input alu;
	input lut;
	input Z;
	input N;
	input C;
	input V;
	output O;
	input CLK;
	input ASYNCRESET;
	wire [0:0] Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst13$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst14$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst15$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst16$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst17$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst18$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst9$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [4:0] const_0_5_out;
	wire [4:0] const_10_5_out;
	wire [4:0] const_11_5_out;
	wire [4:0] const_12_5_out;
	wire [4:0] const_13_5_out;
	wire [4:0] const_14_5_out;
	wire [4:0] const_15_5_out;
	wire [4:0] const_16_5_out;
	wire [4:0] const_17_5_out;
	wire [4:0] const_18_5_out;
	wire [4:0] const_1_5_out;
	wire [4:0] const_2_5_out;
	wire [4:0] const_3_5_out;
	wire [4:0] const_4_5_out;
	wire [4:0] const_5_5_out;
	wire [4:0] const_6_5_out;
	wire [4:0] const_7_5_out;
	wire [4:0] const_8_5_out;
	wire [4:0] const_9_5_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bit_and_inst1_out;
	wire magma_Bit_and_inst2_out;
	wire magma_Bit_and_inst3_out;
	wire magma_Bit_not_inst0_out;
	wire magma_Bit_not_inst1_out;
	wire magma_Bit_not_inst10_out;
	wire magma_Bit_not_inst11_out;
	wire magma_Bit_not_inst12_out;
	wire magma_Bit_not_inst2_out;
	wire magma_Bit_not_inst3_out;
	wire magma_Bit_not_inst4_out;
	wire magma_Bit_not_inst5_out;
	wire magma_Bit_not_inst6_out;
	wire magma_Bit_not_inst7_out;
	wire magma_Bit_not_inst8_out;
	wire magma_Bit_not_inst9_out;
	wire magma_Bit_or_inst0_out;
	wire magma_Bit_or_inst1_out;
	wire magma_Bit_or_inst2_out;
	wire magma_Bit_or_inst3_out;
	wire magma_Bit_or_inst4_out;
	wire magma_Bit_or_inst5_out;
	wire magma_Bit_xor_inst0_out;
	wire magma_Bit_xor_inst1_out;
	wire magma_Bit_xor_inst2_out;
	wire magma_Bit_xor_inst3_out;
	wire magma_Bits_5_eq_inst0_out;
	wire magma_Bits_5_eq_inst1_out;
	wire magma_Bits_5_eq_inst10_out;
	wire magma_Bits_5_eq_inst11_out;
	wire magma_Bits_5_eq_inst12_out;
	wire magma_Bits_5_eq_inst13_out;
	wire magma_Bits_5_eq_inst14_out;
	wire magma_Bits_5_eq_inst15_out;
	wire magma_Bits_5_eq_inst16_out;
	wire magma_Bits_5_eq_inst17_out;
	wire magma_Bits_5_eq_inst18_out;
	wire magma_Bits_5_eq_inst19_out;
	wire magma_Bits_5_eq_inst2_out;
	wire magma_Bits_5_eq_inst20_out;
	wire magma_Bits_5_eq_inst3_out;
	wire magma_Bits_5_eq_inst4_out;
	wire magma_Bits_5_eq_inst5_out;
	wire magma_Bits_5_eq_inst6_out;
	wire magma_Bits_5_eq_inst7_out;
	wire magma_Bits_5_eq_inst8_out;
	wire magma_Bits_5_eq_inst9_out;
	coreir_mux #(.width(1)) Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(magma_Bit_and_inst3_out),
		.in1(magma_Bit_or_inst5_out),
		.sel(magma_Bits_5_eq_inst20_out),
		.out(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(magma_Bit_and_inst2_out),
		.sel(magma_Bits_5_eq_inst19_out),
		.out(Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst10$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst9$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(magma_Bit_and_inst0_out),
		.sel(magma_Bits_5_eq_inst10_out),
		.out(Mux2xBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst11$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(magma_Bit_not_inst3_out),
		.sel(magma_Bits_5_eq_inst9_out),
		.out(Mux2xBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst12$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(V),
		.sel(magma_Bits_5_eq_inst8_out),
		.out(Mux2xBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst13$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(magma_Bit_not_inst2_out),
		.sel(magma_Bits_5_eq_inst7_out),
		.out(Mux2xBit_inst13$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst14$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst13$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(N),
		.sel(magma_Bits_5_eq_inst6_out),
		.out(Mux2xBit_inst14$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst15$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst14$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(magma_Bit_not_inst1_out),
		.sel(magma_Bit_or_inst1_out),
		.out(Mux2xBit_inst15$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst16$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst15$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(C),
		.sel(magma_Bit_or_inst0_out),
		.out(Mux2xBit_inst16$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst17$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst16$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(magma_Bit_not_inst0_out),
		.sel(magma_Bits_5_eq_inst1_out),
		.out(Mux2xBit_inst17$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst18$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst17$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(Z),
		.sel(magma_Bits_5_eq_inst0_out),
		.out(Mux2xBit_inst18$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(magma_Bit_or_inst4_out),
		.sel(magma_Bits_5_eq_inst18_out),
		.out(Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(lut),
		.sel(magma_Bits_5_eq_inst17_out),
		.out(Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(alu),
		.sel(magma_Bits_5_eq_inst16_out),
		.out(Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst5$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(magma_Bit_or_inst3_out),
		.sel(magma_Bits_5_eq_inst15_out),
		.out(Mux2xBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst6$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(magma_Bit_and_inst1_out),
		.sel(magma_Bits_5_eq_inst14_out),
		.out(Mux2xBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst7$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(magma_Bit_xor_inst1_out),
		.sel(magma_Bits_5_eq_inst13_out),
		.out(Mux2xBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst8$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(magma_Bit_not_inst6_out),
		.sel(magma_Bits_5_eq_inst12_out),
		.out(Mux2xBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst9$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(magma_Bit_or_inst2_out),
		.sel(magma_Bits_5_eq_inst11_out),
		.out(Mux2xBit_inst9$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_const #(
		.value(5'h00),
		.width(5)
	) const_0_5(.out(const_0_5_out));
	coreir_const #(
		.value(5'h0a),
		.width(5)
	) const_10_5(.out(const_10_5_out));
	coreir_const #(
		.value(5'h0b),
		.width(5)
	) const_11_5(.out(const_11_5_out));
	coreir_const #(
		.value(5'h0c),
		.width(5)
	) const_12_5(.out(const_12_5_out));
	coreir_const #(
		.value(5'h0d),
		.width(5)
	) const_13_5(.out(const_13_5_out));
	coreir_const #(
		.value(5'h0e),
		.width(5)
	) const_14_5(.out(const_14_5_out));
	coreir_const #(
		.value(5'h0f),
		.width(5)
	) const_15_5(.out(const_15_5_out));
	coreir_const #(
		.value(5'h10),
		.width(5)
	) const_16_5(.out(const_16_5_out));
	coreir_const #(
		.value(5'h11),
		.width(5)
	) const_17_5(.out(const_17_5_out));
	coreir_const #(
		.value(5'h12),
		.width(5)
	) const_18_5(.out(const_18_5_out));
	coreir_const #(
		.value(5'h01),
		.width(5)
	) const_1_5(.out(const_1_5_out));
	coreir_const #(
		.value(5'h02),
		.width(5)
	) const_2_5(.out(const_2_5_out));
	coreir_const #(
		.value(5'h03),
		.width(5)
	) const_3_5(.out(const_3_5_out));
	coreir_const #(
		.value(5'h04),
		.width(5)
	) const_4_5(.out(const_4_5_out));
	coreir_const #(
		.value(5'h05),
		.width(5)
	) const_5_5(.out(const_5_5_out));
	coreir_const #(
		.value(5'h06),
		.width(5)
	) const_6_5(.out(const_6_5_out));
	coreir_const #(
		.value(5'h07),
		.width(5)
	) const_7_5(.out(const_7_5_out));
	coreir_const #(
		.value(5'h08),
		.width(5)
	) const_8_5(.out(const_8_5_out));
	coreir_const #(
		.value(5'h09),
		.width(5)
	) const_9_5(.out(const_9_5_out));
	corebit_and magma_Bit_and_inst0(
		.in0(C),
		.in1(magma_Bit_not_inst4_out),
		.out(magma_Bit_and_inst0_out)
	);
	corebit_and magma_Bit_and_inst1(
		.in0(magma_Bit_not_inst7_out),
		.in1(magma_Bit_not_inst8_out),
		.out(magma_Bit_and_inst1_out)
	);
	corebit_and magma_Bit_and_inst2(
		.in0(magma_Bit_not_inst10_out),
		.in1(magma_Bit_not_inst11_out),
		.out(magma_Bit_and_inst2_out)
	);
	corebit_and magma_Bit_and_inst3(
		.in0(N),
		.in1(magma_Bit_not_inst12_out),
		.out(magma_Bit_and_inst3_out)
	);
	corebit_not magma_Bit_not_inst0(
		.in(Z),
		.out(magma_Bit_not_inst0_out)
	);
	corebit_not magma_Bit_not_inst1(
		.in(C),
		.out(magma_Bit_not_inst1_out)
	);
	corebit_not magma_Bit_not_inst10(
		.in(N),
		.out(magma_Bit_not_inst10_out)
	);
	corebit_not magma_Bit_not_inst11(
		.in(Z),
		.out(magma_Bit_not_inst11_out)
	);
	corebit_not magma_Bit_not_inst12(
		.in(Z),
		.out(magma_Bit_not_inst12_out)
	);
	corebit_not magma_Bit_not_inst2(
		.in(N),
		.out(magma_Bit_not_inst2_out)
	);
	corebit_not magma_Bit_not_inst3(
		.in(V),
		.out(magma_Bit_not_inst3_out)
	);
	corebit_not magma_Bit_not_inst4(
		.in(Z),
		.out(magma_Bit_not_inst4_out)
	);
	corebit_not magma_Bit_not_inst5(
		.in(C),
		.out(magma_Bit_not_inst5_out)
	);
	corebit_not magma_Bit_not_inst6(
		.in(magma_Bit_xor_inst0_out),
		.out(magma_Bit_not_inst6_out)
	);
	corebit_not magma_Bit_not_inst7(
		.in(Z),
		.out(magma_Bit_not_inst7_out)
	);
	corebit_not magma_Bit_not_inst8(
		.in(magma_Bit_xor_inst2_out),
		.out(magma_Bit_not_inst8_out)
	);
	corebit_not magma_Bit_not_inst9(
		.in(N),
		.out(magma_Bit_not_inst9_out)
	);
	corebit_or magma_Bit_or_inst0(
		.in0(magma_Bits_5_eq_inst2_out),
		.in1(magma_Bits_5_eq_inst3_out),
		.out(magma_Bit_or_inst0_out)
	);
	corebit_or magma_Bit_or_inst1(
		.in0(magma_Bits_5_eq_inst4_out),
		.in1(magma_Bits_5_eq_inst5_out),
		.out(magma_Bit_or_inst1_out)
	);
	corebit_or magma_Bit_or_inst2(
		.in0(magma_Bit_not_inst5_out),
		.in1(Z),
		.out(magma_Bit_or_inst2_out)
	);
	corebit_or magma_Bit_or_inst3(
		.in0(Z),
		.in1(magma_Bit_xor_inst3_out),
		.out(magma_Bit_or_inst3_out)
	);
	corebit_or magma_Bit_or_inst4(
		.in0(magma_Bit_not_inst9_out),
		.in1(Z),
		.out(magma_Bit_or_inst4_out)
	);
	corebit_or magma_Bit_or_inst5(
		.in0(N),
		.in1(Z),
		.out(magma_Bit_or_inst5_out)
	);
	corebit_xor magma_Bit_xor_inst0(
		.in0(N),
		.in1(V),
		.out(magma_Bit_xor_inst0_out)
	);
	corebit_xor magma_Bit_xor_inst1(
		.in0(N),
		.in1(V),
		.out(magma_Bit_xor_inst1_out)
	);
	corebit_xor magma_Bit_xor_inst2(
		.in0(N),
		.in1(V),
		.out(magma_Bit_xor_inst2_out)
	);
	corebit_xor magma_Bit_xor_inst3(
		.in0(N),
		.in1(V),
		.out(magma_Bit_xor_inst3_out)
	);
	coreir_eq #(.width(5)) magma_Bits_5_eq_inst0(
		.in0(code),
		.in1(const_0_5_out),
		.out(magma_Bits_5_eq_inst0_out)
	);
	coreir_eq #(.width(5)) magma_Bits_5_eq_inst1(
		.in0(code),
		.in1(const_1_5_out),
		.out(magma_Bits_5_eq_inst1_out)
	);
	coreir_eq #(.width(5)) magma_Bits_5_eq_inst10(
		.in0(code),
		.in1(const_8_5_out),
		.out(magma_Bits_5_eq_inst10_out)
	);
	coreir_eq #(.width(5)) magma_Bits_5_eq_inst11(
		.in0(code),
		.in1(const_9_5_out),
		.out(magma_Bits_5_eq_inst11_out)
	);
	coreir_eq #(.width(5)) magma_Bits_5_eq_inst12(
		.in0(code),
		.in1(const_10_5_out),
		.out(magma_Bits_5_eq_inst12_out)
	);
	coreir_eq #(.width(5)) magma_Bits_5_eq_inst13(
		.in0(code),
		.in1(const_11_5_out),
		.out(magma_Bits_5_eq_inst13_out)
	);
	coreir_eq #(.width(5)) magma_Bits_5_eq_inst14(
		.in0(code),
		.in1(const_12_5_out),
		.out(magma_Bits_5_eq_inst14_out)
	);
	coreir_eq #(.width(5)) magma_Bits_5_eq_inst15(
		.in0(code),
		.in1(const_13_5_out),
		.out(magma_Bits_5_eq_inst15_out)
	);
	coreir_eq #(.width(5)) magma_Bits_5_eq_inst16(
		.in0(code),
		.in1(const_15_5_out),
		.out(magma_Bits_5_eq_inst16_out)
	);
	coreir_eq #(.width(5)) magma_Bits_5_eq_inst17(
		.in0(code),
		.in1(const_14_5_out),
		.out(magma_Bits_5_eq_inst17_out)
	);
	coreir_eq #(.width(5)) magma_Bits_5_eq_inst18(
		.in0(code),
		.in1(const_16_5_out),
		.out(magma_Bits_5_eq_inst18_out)
	);
	coreir_eq #(.width(5)) magma_Bits_5_eq_inst19(
		.in0(code),
		.in1(const_17_5_out),
		.out(magma_Bits_5_eq_inst19_out)
	);
	coreir_eq #(.width(5)) magma_Bits_5_eq_inst2(
		.in0(code),
		.in1(const_2_5_out),
		.out(magma_Bits_5_eq_inst2_out)
	);
	coreir_eq #(.width(5)) magma_Bits_5_eq_inst20(
		.in0(code),
		.in1(const_18_5_out),
		.out(magma_Bits_5_eq_inst20_out)
	);
	coreir_eq #(.width(5)) magma_Bits_5_eq_inst3(
		.in0(code),
		.in1(const_2_5_out),
		.out(magma_Bits_5_eq_inst3_out)
	);
	coreir_eq #(.width(5)) magma_Bits_5_eq_inst4(
		.in0(code),
		.in1(const_3_5_out),
		.out(magma_Bits_5_eq_inst4_out)
	);
	coreir_eq #(.width(5)) magma_Bits_5_eq_inst5(
		.in0(code),
		.in1(const_3_5_out),
		.out(magma_Bits_5_eq_inst5_out)
	);
	coreir_eq #(.width(5)) magma_Bits_5_eq_inst6(
		.in0(code),
		.in1(const_4_5_out),
		.out(magma_Bits_5_eq_inst6_out)
	);
	coreir_eq #(.width(5)) magma_Bits_5_eq_inst7(
		.in0(code),
		.in1(const_5_5_out),
		.out(magma_Bits_5_eq_inst7_out)
	);
	coreir_eq #(.width(5)) magma_Bits_5_eq_inst8(
		.in0(code),
		.in1(const_6_5_out),
		.out(magma_Bits_5_eq_inst8_out)
	);
	coreir_eq #(.width(5)) magma_Bits_5_eq_inst9(
		.in0(code),
		.in1(const_7_5_out),
		.out(magma_Bits_5_eq_inst9_out)
	);
	assign O = Mux2xBit_inst18$coreir_commonlib_mux2x1_inst0$_join_out[0];
endmodule
module CB_input_width_1_num_1_sel (
	I,
	O
);
	input [3:0] I;
	output [3:0] O;
	assign O = I;
endmodule
module CB_input_width_1_num_1 (
	I_0,
	I_1,
	I_10,
	I_11,
	I_2,
	I_3,
	I_4,
	I_5,
	I_6,
	I_7,
	I_8,
	I_9,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	read_config_data,
	reset
);
	input [0:0] I_0;
	input [0:0] I_1;
	input [0:0] I_10;
	input [0:0] I_11;
	input [0:0] I_2;
	input [0:0] I_3;
	input [0:0] I_4;
	input [0:0] I_5;
	input [0:0] I_6;
	input [0:0] I_7;
	input [0:0] I_8;
	input [0:0] I_9;
	output [0:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output [31:0] read_config_data;
	input reset;
	wire [3:0] CB_input_width_1_num_1_sel_inst0_O;
	wire [0:0] MUX_CB_input_width_1_num_1$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0_out;
	wire ZextWrapper_4_32_inst0$bit_const_0_None_out;
	wire [3:0] ZextWrapper_4_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_4_32_inst0$self_O_in;
	wire [3:0] config_reg_0_O;
	CB_input_width_1_num_1_sel CB_input_width_1_num_1_sel_inst0(
		.I(config_reg_0_O),
		.O(CB_input_width_1_num_1_sel_inst0_O)
	);
	commonlib_muxn__N12__width1 MUX_CB_input_width_1_num_1$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0(
		.in_data_0(I_0),
		.in_data_1(I_1),
		.in_data_10(I_10),
		.in_data_11(I_11),
		.in_data_2(I_2),
		.in_data_3(I_3),
		.in_data_4(I_4),
		.in_data_5(I_5),
		.in_data_6(I_6),
		.in_data_7(I_7),
		.in_data_8(I_8),
		.in_data_9(I_9),
		.in_sel(CB_input_width_1_num_1_sel_inst0_O),
		.out(MUX_CB_input_width_1_num_1$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_4_32_inst0$bit_const_0_None(.out(ZextWrapper_4_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit4 ZextWrapper_4_32_inst0$self_I(
		.in(config_reg_0_O),
		.out(ZextWrapper_4_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_4_32_inst0$self_O_out;
	assign ZextWrapper_4_32_inst0$self_O_out = {ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$self_I_out[3:0]};
	mantle_wire__typeBitIn32 ZextWrapper_4_32_inst0$self_O(
		.in(ZextWrapper_4_32_inst0$self_O_in),
		.out(ZextWrapper_4_32_inst0$self_O_out)
	);
	ConfigRegister_4_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = MUX_CB_input_width_1_num_1$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0_out;
	assign read_config_data = ZextWrapper_4_32_inst0$self_O_in;
endmodule
module CB_input_width_1_num_0_sel (
	I,
	O
);
	input [3:0] I;
	output [3:0] O;
	assign O = I;
endmodule
module CB_input_width_1_num_0 (
	I_0,
	I_1,
	I_10,
	I_11,
	I_2,
	I_3,
	I_4,
	I_5,
	I_6,
	I_7,
	I_8,
	I_9,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	read_config_data,
	reset
);
	input [0:0] I_0;
	input [0:0] I_1;
	input [0:0] I_10;
	input [0:0] I_11;
	input [0:0] I_2;
	input [0:0] I_3;
	input [0:0] I_4;
	input [0:0] I_5;
	input [0:0] I_6;
	input [0:0] I_7;
	input [0:0] I_8;
	input [0:0] I_9;
	output [0:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output [31:0] read_config_data;
	input reset;
	wire [3:0] CB_input_width_1_num_0_sel_inst0_O;
	wire [0:0] MUX_CB_input_width_1_num_0$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0_out;
	wire ZextWrapper_4_32_inst0$bit_const_0_None_out;
	wire [3:0] ZextWrapper_4_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_4_32_inst0$self_O_in;
	wire [3:0] config_reg_0_O;
	CB_input_width_1_num_0_sel CB_input_width_1_num_0_sel_inst0(
		.I(config_reg_0_O),
		.O(CB_input_width_1_num_0_sel_inst0_O)
	);
	commonlib_muxn__N12__width1 MUX_CB_input_width_1_num_0$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0(
		.in_data_0(I_0),
		.in_data_1(I_1),
		.in_data_10(I_10),
		.in_data_11(I_11),
		.in_data_2(I_2),
		.in_data_3(I_3),
		.in_data_4(I_4),
		.in_data_5(I_5),
		.in_data_6(I_6),
		.in_data_7(I_7),
		.in_data_8(I_8),
		.in_data_9(I_9),
		.in_sel(CB_input_width_1_num_0_sel_inst0_O),
		.out(MUX_CB_input_width_1_num_0$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_4_32_inst0$bit_const_0_None(.out(ZextWrapper_4_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit4 ZextWrapper_4_32_inst0$self_I(
		.in(config_reg_0_O),
		.out(ZextWrapper_4_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_4_32_inst0$self_O_out;
	assign ZextWrapper_4_32_inst0$self_O_out = {ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$self_I_out[3:0]};
	mantle_wire__typeBitIn32 ZextWrapper_4_32_inst0$self_O(
		.in(ZextWrapper_4_32_inst0$self_O_in),
		.out(ZextWrapper_4_32_inst0$self_O_out)
	);
	ConfigRegister_4_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = MUX_CB_input_width_1_num_0$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0_out;
	assign read_config_data = ZextWrapper_4_32_inst0$self_O_in;
endmodule
module CB_input_width_16_num_3_sel (
	I,
	O
);
	input [3:0] I;
	output [3:0] O;
	assign O = I;
endmodule
module CB_input_width_16_num_3 (
	I_0,
	I_1,
	I_10,
	I_11,
	I_2,
	I_3,
	I_4,
	I_5,
	I_6,
	I_7,
	I_8,
	I_9,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	read_config_data,
	reset
);
	input [15:0] I_0;
	input [15:0] I_1;
	input [15:0] I_10;
	input [15:0] I_11;
	input [15:0] I_2;
	input [15:0] I_3;
	input [15:0] I_4;
	input [15:0] I_5;
	input [15:0] I_6;
	input [15:0] I_7;
	input [15:0] I_8;
	input [15:0] I_9;
	output [15:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output [31:0] read_config_data;
	input reset;
	wire [3:0] CB_input_width_16_num_3_sel_inst0_O;
	wire [15:0] MUX_CB_input_width_16_num_3$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0_out;
	wire ZextWrapper_4_32_inst0$bit_const_0_None_out;
	wire [3:0] ZextWrapper_4_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_4_32_inst0$self_O_in;
	wire [3:0] config_reg_0_O;
	CB_input_width_16_num_3_sel CB_input_width_16_num_3_sel_inst0(
		.I(config_reg_0_O),
		.O(CB_input_width_16_num_3_sel_inst0_O)
	);
	commonlib_muxn__N12__width16 MUX_CB_input_width_16_num_3$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0(
		.in_data_0(I_0),
		.in_data_1(I_1),
		.in_data_10(I_10),
		.in_data_11(I_11),
		.in_data_2(I_2),
		.in_data_3(I_3),
		.in_data_4(I_4),
		.in_data_5(I_5),
		.in_data_6(I_6),
		.in_data_7(I_7),
		.in_data_8(I_8),
		.in_data_9(I_9),
		.in_sel(CB_input_width_16_num_3_sel_inst0_O),
		.out(MUX_CB_input_width_16_num_3$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_4_32_inst0$bit_const_0_None(.out(ZextWrapper_4_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit4 ZextWrapper_4_32_inst0$self_I(
		.in(config_reg_0_O),
		.out(ZextWrapper_4_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_4_32_inst0$self_O_out;
	assign ZextWrapper_4_32_inst0$self_O_out = {ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$self_I_out[3:0]};
	mantle_wire__typeBitIn32 ZextWrapper_4_32_inst0$self_O(
		.in(ZextWrapper_4_32_inst0$self_O_in),
		.out(ZextWrapper_4_32_inst0$self_O_out)
	);
	ConfigRegister_4_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = MUX_CB_input_width_16_num_3$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0_out;
	assign read_config_data = ZextWrapper_4_32_inst0$self_O_in;
endmodule
module CB_input_width_16_num_2_sel (
	I,
	O
);
	input [3:0] I;
	output [3:0] O;
	assign O = I;
endmodule
module CB_input_width_16_num_2 (
	I_0,
	I_1,
	I_10,
	I_11,
	I_2,
	I_3,
	I_4,
	I_5,
	I_6,
	I_7,
	I_8,
	I_9,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	read_config_data,
	reset
);
	input [15:0] I_0;
	input [15:0] I_1;
	input [15:0] I_10;
	input [15:0] I_11;
	input [15:0] I_2;
	input [15:0] I_3;
	input [15:0] I_4;
	input [15:0] I_5;
	input [15:0] I_6;
	input [15:0] I_7;
	input [15:0] I_8;
	input [15:0] I_9;
	output [15:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output [31:0] read_config_data;
	input reset;
	wire [3:0] CB_input_width_16_num_2_sel_inst0_O;
	wire [15:0] MUX_CB_input_width_16_num_2$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0_out;
	wire ZextWrapper_4_32_inst0$bit_const_0_None_out;
	wire [3:0] ZextWrapper_4_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_4_32_inst0$self_O_in;
	wire [3:0] config_reg_0_O;
	CB_input_width_16_num_2_sel CB_input_width_16_num_2_sel_inst0(
		.I(config_reg_0_O),
		.O(CB_input_width_16_num_2_sel_inst0_O)
	);
	commonlib_muxn__N12__width16 MUX_CB_input_width_16_num_2$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0(
		.in_data_0(I_0),
		.in_data_1(I_1),
		.in_data_10(I_10),
		.in_data_11(I_11),
		.in_data_2(I_2),
		.in_data_3(I_3),
		.in_data_4(I_4),
		.in_data_5(I_5),
		.in_data_6(I_6),
		.in_data_7(I_7),
		.in_data_8(I_8),
		.in_data_9(I_9),
		.in_sel(CB_input_width_16_num_2_sel_inst0_O),
		.out(MUX_CB_input_width_16_num_2$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_4_32_inst0$bit_const_0_None(.out(ZextWrapper_4_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit4 ZextWrapper_4_32_inst0$self_I(
		.in(config_reg_0_O),
		.out(ZextWrapper_4_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_4_32_inst0$self_O_out;
	assign ZextWrapper_4_32_inst0$self_O_out = {ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$self_I_out[3:0]};
	mantle_wire__typeBitIn32 ZextWrapper_4_32_inst0$self_O(
		.in(ZextWrapper_4_32_inst0$self_O_in),
		.out(ZextWrapper_4_32_inst0$self_O_out)
	);
	ConfigRegister_4_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = MUX_CB_input_width_16_num_2$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0_out;
	assign read_config_data = ZextWrapper_4_32_inst0$self_O_in;
endmodule
module CB_input_width_16_num_1_sel (
	I,
	O
);
	input [3:0] I;
	output [3:0] O;
	assign O = I;
endmodule
module CB_input_width_16_num_1 (
	I_0,
	I_1,
	I_10,
	I_11,
	I_2,
	I_3,
	I_4,
	I_5,
	I_6,
	I_7,
	I_8,
	I_9,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	read_config_data,
	reset
);
	input [15:0] I_0;
	input [15:0] I_1;
	input [15:0] I_10;
	input [15:0] I_11;
	input [15:0] I_2;
	input [15:0] I_3;
	input [15:0] I_4;
	input [15:0] I_5;
	input [15:0] I_6;
	input [15:0] I_7;
	input [15:0] I_8;
	input [15:0] I_9;
	output [15:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output [31:0] read_config_data;
	input reset;
	wire [3:0] CB_input_width_16_num_1_sel_inst0_O;
	wire [15:0] MUX_CB_input_width_16_num_1$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0_out;
	wire ZextWrapper_4_32_inst0$bit_const_0_None_out;
	wire [3:0] ZextWrapper_4_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_4_32_inst0$self_O_in;
	wire [3:0] config_reg_0_O;
	CB_input_width_16_num_1_sel CB_input_width_16_num_1_sel_inst0(
		.I(config_reg_0_O),
		.O(CB_input_width_16_num_1_sel_inst0_O)
	);
	commonlib_muxn__N12__width16 MUX_CB_input_width_16_num_1$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0(
		.in_data_0(I_0),
		.in_data_1(I_1),
		.in_data_10(I_10),
		.in_data_11(I_11),
		.in_data_2(I_2),
		.in_data_3(I_3),
		.in_data_4(I_4),
		.in_data_5(I_5),
		.in_data_6(I_6),
		.in_data_7(I_7),
		.in_data_8(I_8),
		.in_data_9(I_9),
		.in_sel(CB_input_width_16_num_1_sel_inst0_O),
		.out(MUX_CB_input_width_16_num_1$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_4_32_inst0$bit_const_0_None(.out(ZextWrapper_4_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit4 ZextWrapper_4_32_inst0$self_I(
		.in(config_reg_0_O),
		.out(ZextWrapper_4_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_4_32_inst0$self_O_out;
	assign ZextWrapper_4_32_inst0$self_O_out = {ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$self_I_out[3:0]};
	mantle_wire__typeBitIn32 ZextWrapper_4_32_inst0$self_O(
		.in(ZextWrapper_4_32_inst0$self_O_in),
		.out(ZextWrapper_4_32_inst0$self_O_out)
	);
	ConfigRegister_4_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = MUX_CB_input_width_16_num_1$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0_out;
	assign read_config_data = ZextWrapper_4_32_inst0$self_O_in;
endmodule
module CB_input_width_16_num_0_sel (
	I,
	O
);
	input [3:0] I;
	output [3:0] O;
	assign O = I;
endmodule
module CB_input_width_16_num_0 (
	I_0,
	I_1,
	I_10,
	I_11,
	I_2,
	I_3,
	I_4,
	I_5,
	I_6,
	I_7,
	I_8,
	I_9,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	read_config_data,
	reset
);
	input [15:0] I_0;
	input [15:0] I_1;
	input [15:0] I_10;
	input [15:0] I_11;
	input [15:0] I_2;
	input [15:0] I_3;
	input [15:0] I_4;
	input [15:0] I_5;
	input [15:0] I_6;
	input [15:0] I_7;
	input [15:0] I_8;
	input [15:0] I_9;
	output [15:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output [31:0] read_config_data;
	input reset;
	wire [3:0] CB_input_width_16_num_0_sel_inst0_O;
	wire [15:0] MUX_CB_input_width_16_num_0$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0_out;
	wire ZextWrapper_4_32_inst0$bit_const_0_None_out;
	wire [3:0] ZextWrapper_4_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_4_32_inst0$self_O_in;
	wire [3:0] config_reg_0_O;
	CB_input_width_16_num_0_sel CB_input_width_16_num_0_sel_inst0(
		.I(config_reg_0_O),
		.O(CB_input_width_16_num_0_sel_inst0_O)
	);
	commonlib_muxn__N12__width16 MUX_CB_input_width_16_num_0$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0(
		.in_data_0(I_0),
		.in_data_1(I_1),
		.in_data_10(I_10),
		.in_data_11(I_11),
		.in_data_2(I_2),
		.in_data_3(I_3),
		.in_data_4(I_4),
		.in_data_5(I_5),
		.in_data_6(I_6),
		.in_data_7(I_7),
		.in_data_8(I_8),
		.in_data_9(I_9),
		.in_sel(CB_input_width_16_num_0_sel_inst0_O),
		.out(MUX_CB_input_width_16_num_0$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_4_32_inst0$bit_const_0_None(.out(ZextWrapper_4_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit4 ZextWrapper_4_32_inst0$self_I(
		.in(config_reg_0_O),
		.out(ZextWrapper_4_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_4_32_inst0$self_O_out;
	assign ZextWrapper_4_32_inst0$self_O_out = {ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$self_I_out[3:0]};
	mantle_wire__typeBitIn32 ZextWrapper_4_32_inst0$self_O(
		.in(ZextWrapper_4_32_inst0$self_O_in),
		.out(ZextWrapper_4_32_inst0$self_O_out)
	);
	ConfigRegister_4_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = MUX_CB_input_width_16_num_0$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0_out;
	assign read_config_data = ZextWrapper_4_32_inst0$self_O_in;
endmodule
module CB_flush_sel (
	I,
	O
);
	input [3:0] I;
	output [3:0] O;
	assign O = I;
endmodule
module CB_flush (
	I_0,
	I_1,
	I_10,
	I_11,
	I_2,
	I_3,
	I_4,
	I_5,
	I_6,
	I_7,
	I_8,
	I_9,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	read_config_data,
	reset
);
	input [0:0] I_0;
	input [0:0] I_1;
	input [0:0] I_10;
	input [0:0] I_11;
	input [0:0] I_2;
	input [0:0] I_3;
	input [0:0] I_4;
	input [0:0] I_5;
	input [0:0] I_6;
	input [0:0] I_7;
	input [0:0] I_8;
	input [0:0] I_9;
	output [0:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output [31:0] read_config_data;
	input reset;
	wire [3:0] CB_flush_sel_inst0_O;
	wire [0:0] MUX_CB_flush$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0_out;
	wire ZextWrapper_4_32_inst0$bit_const_0_None_out;
	wire [3:0] ZextWrapper_4_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_4_32_inst0$self_O_in;
	wire [3:0] config_reg_0_O;
	CB_flush_sel CB_flush_sel_inst0(
		.I(config_reg_0_O),
		.O(CB_flush_sel_inst0_O)
	);
	commonlib_muxn__N12__width1 MUX_CB_flush$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0(
		.in_data_0(I_0),
		.in_data_1(I_1),
		.in_data_10(I_10),
		.in_data_11(I_11),
		.in_data_2(I_2),
		.in_data_3(I_3),
		.in_data_4(I_4),
		.in_data_5(I_5),
		.in_data_6(I_6),
		.in_data_7(I_7),
		.in_data_8(I_8),
		.in_data_9(I_9),
		.in_sel(CB_flush_sel_inst0_O),
		.out(MUX_CB_flush$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_4_32_inst0$bit_const_0_None(.out(ZextWrapper_4_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit4 ZextWrapper_4_32_inst0$self_I(
		.in(config_reg_0_O),
		.out(ZextWrapper_4_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_4_32_inst0$self_O_out;
	assign ZextWrapper_4_32_inst0$self_O_out = {ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$self_I_out[3:0]};
	mantle_wire__typeBitIn32 ZextWrapper_4_32_inst0$self_O(
		.in(ZextWrapper_4_32_inst0$self_O_in),
		.out(ZextWrapper_4_32_inst0$self_O_out)
	);
	ConfigRegister_4_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = MUX_CB_flush$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0_out;
	assign read_config_data = ZextWrapper_4_32_inst0$self_O_in;
endmodule
module Tile_MemCore (
	SB_T0_EAST_SB_IN_B1,
	SB_T0_EAST_SB_IN_B16,
	SB_T0_EAST_SB_OUT_B1,
	SB_T0_EAST_SB_OUT_B16,
	SB_T0_NORTH_SB_IN_B1,
	SB_T0_NORTH_SB_IN_B16,
	SB_T0_NORTH_SB_OUT_B1,
	SB_T0_NORTH_SB_OUT_B16,
	SB_T0_SOUTH_SB_IN_B1,
	SB_T0_SOUTH_SB_IN_B16,
	SB_T0_SOUTH_SB_OUT_B1,
	SB_T0_SOUTH_SB_OUT_B16,
	SB_T0_WEST_SB_IN_B1,
	SB_T0_WEST_SB_IN_B16,
	SB_T0_WEST_SB_OUT_B1,
	SB_T0_WEST_SB_OUT_B16,
	SB_T1_EAST_SB_IN_B1,
	SB_T1_EAST_SB_IN_B16,
	SB_T1_EAST_SB_OUT_B1,
	SB_T1_EAST_SB_OUT_B16,
	SB_T1_NORTH_SB_IN_B1,
	SB_T1_NORTH_SB_IN_B16,
	SB_T1_NORTH_SB_OUT_B1,
	SB_T1_NORTH_SB_OUT_B16,
	SB_T1_SOUTH_SB_IN_B1,
	SB_T1_SOUTH_SB_IN_B16,
	SB_T1_SOUTH_SB_OUT_B1,
	SB_T1_SOUTH_SB_OUT_B16,
	SB_T1_WEST_SB_IN_B1,
	SB_T1_WEST_SB_IN_B16,
	SB_T1_WEST_SB_OUT_B1,
	SB_T1_WEST_SB_OUT_B16,
	SB_T2_EAST_SB_IN_B1,
	SB_T2_EAST_SB_IN_B16,
	SB_T2_EAST_SB_OUT_B1,
	SB_T2_EAST_SB_OUT_B16,
	SB_T2_NORTH_SB_IN_B1,
	SB_T2_NORTH_SB_IN_B16,
	SB_T2_NORTH_SB_OUT_B1,
	SB_T2_NORTH_SB_OUT_B16,
	SB_T2_SOUTH_SB_IN_B1,
	SB_T2_SOUTH_SB_IN_B16,
	SB_T2_SOUTH_SB_OUT_B1,
	SB_T2_SOUTH_SB_OUT_B16,
	SB_T2_WEST_SB_IN_B1,
	SB_T2_WEST_SB_IN_B16,
	SB_T2_WEST_SB_OUT_B1,
	SB_T2_WEST_SB_OUT_B16,
	clk,
	clk_out,
	clk_pass_through,
	clk_pass_through_out_bot,
	config_config_addr,
	config_config_data,
	config_out_config_addr,
	config_out_config_data,
	config_out_read,
	config_out_write,
	config_read,
	config_write,
	hi,
	lo,
	read_config_data,
	read_config_data_in,
	reset,
	reset_out,
	stall,
	stall_out,
	tile_id
);
	input [0:0] SB_T0_EAST_SB_IN_B1;
	input [15:0] SB_T0_EAST_SB_IN_B16;
	output [0:0] SB_T0_EAST_SB_OUT_B1;
	output [15:0] SB_T0_EAST_SB_OUT_B16;
	input [0:0] SB_T0_NORTH_SB_IN_B1;
	input [15:0] SB_T0_NORTH_SB_IN_B16;
	output [0:0] SB_T0_NORTH_SB_OUT_B1;
	output [15:0] SB_T0_NORTH_SB_OUT_B16;
	input [0:0] SB_T0_SOUTH_SB_IN_B1;
	input [15:0] SB_T0_SOUTH_SB_IN_B16;
	output [0:0] SB_T0_SOUTH_SB_OUT_B1;
	output [15:0] SB_T0_SOUTH_SB_OUT_B16;
	input [0:0] SB_T0_WEST_SB_IN_B1;
	input [15:0] SB_T0_WEST_SB_IN_B16;
	output [0:0] SB_T0_WEST_SB_OUT_B1;
	output [15:0] SB_T0_WEST_SB_OUT_B16;
	input [0:0] SB_T1_EAST_SB_IN_B1;
	input [15:0] SB_T1_EAST_SB_IN_B16;
	output [0:0] SB_T1_EAST_SB_OUT_B1;
	output [15:0] SB_T1_EAST_SB_OUT_B16;
	input [0:0] SB_T1_NORTH_SB_IN_B1;
	input [15:0] SB_T1_NORTH_SB_IN_B16;
	output [0:0] SB_T1_NORTH_SB_OUT_B1;
	output [15:0] SB_T1_NORTH_SB_OUT_B16;
	input [0:0] SB_T1_SOUTH_SB_IN_B1;
	input [15:0] SB_T1_SOUTH_SB_IN_B16;
	output [0:0] SB_T1_SOUTH_SB_OUT_B1;
	output [15:0] SB_T1_SOUTH_SB_OUT_B16;
	input [0:0] SB_T1_WEST_SB_IN_B1;
	input [15:0] SB_T1_WEST_SB_IN_B16;
	output [0:0] SB_T1_WEST_SB_OUT_B1;
	output [15:0] SB_T1_WEST_SB_OUT_B16;
	input [0:0] SB_T2_EAST_SB_IN_B1;
	input [15:0] SB_T2_EAST_SB_IN_B16;
	output [0:0] SB_T2_EAST_SB_OUT_B1;
	output [15:0] SB_T2_EAST_SB_OUT_B16;
	input [0:0] SB_T2_NORTH_SB_IN_B1;
	input [15:0] SB_T2_NORTH_SB_IN_B16;
	output [0:0] SB_T2_NORTH_SB_OUT_B1;
	output [15:0] SB_T2_NORTH_SB_OUT_B16;
	input [0:0] SB_T2_SOUTH_SB_IN_B1;
	input [15:0] SB_T2_SOUTH_SB_IN_B16;
	output [0:0] SB_T2_SOUTH_SB_OUT_B1;
	output [15:0] SB_T2_SOUTH_SB_OUT_B16;
	input [0:0] SB_T2_WEST_SB_IN_B1;
	input [15:0] SB_T2_WEST_SB_IN_B16;
	output [0:0] SB_T2_WEST_SB_OUT_B1;
	output [15:0] SB_T2_WEST_SB_OUT_B16;
	input clk;
	output clk_out;
	input clk_pass_through;
	output clk_pass_through_out_bot;
	input [31:0] config_config_addr;
	input [31:0] config_config_data;
	output [31:0] config_out_config_addr;
	output [31:0] config_out_config_data;
	output [0:0] config_out_read;
	output [0:0] config_out_write;
	input [0:0] config_read;
	input [0:0] config_write;
	output [8:0] hi;
	output [7:0] lo;
	output [31:0] read_config_data;
	input [31:0] read_config_data_in;
	input reset;
	output reset_out;
	input [0:0] stall;
	output [0:0] stall_out;
	input [15:0] tile_id;
	wire [0:0] CB_flush_O;
	wire [31:0] CB_flush_read_config_data;
	wire [7:0] CB_flush_config_config_addr_in;
	wire [15:0] CB_input_width_16_num_0_O;
	wire [31:0] CB_input_width_16_num_0_read_config_data;
	wire [7:0] CB_input_width_16_num_0_config_config_addr_in;
	wire [15:0] CB_input_width_16_num_1_O;
	wire [31:0] CB_input_width_16_num_1_read_config_data;
	wire [7:0] CB_input_width_16_num_1_config_config_addr_in;
	wire [15:0] CB_input_width_16_num_2_O;
	wire [31:0] CB_input_width_16_num_2_read_config_data;
	wire [7:0] CB_input_width_16_num_2_config_config_addr_in;
	wire [15:0] CB_input_width_16_num_3_O;
	wire [31:0] CB_input_width_16_num_3_read_config_data;
	wire [7:0] CB_input_width_16_num_3_config_config_addr_in;
	wire [0:0] CB_input_width_1_num_0_O;
	wire [31:0] CB_input_width_1_num_0_read_config_data;
	wire [7:0] CB_input_width_1_num_0_config_config_addr_in;
	wire [0:0] CB_input_width_1_num_1_O;
	wire [31:0] CB_input_width_1_num_1_read_config_data;
	wire [7:0] CB_input_width_1_num_1_config_config_addr_in;
	wire DECODE_FEATURE_0_O;
	wire DECODE_FEATURE_1_O;
	wire DECODE_FEATURE_10_O;
	wire DECODE_FEATURE_2_O;
	wire DECODE_FEATURE_3_O;
	wire DECODE_FEATURE_4_O;
	wire DECODE_FEATURE_5_O;
	wire DECODE_FEATURE_6_O;
	wire DECODE_FEATURE_7_O;
	wire DECODE_FEATURE_8_O;
	wire DECODE_FEATURE_9_O;
	wire FEATURE_AND_0_out;
	wire FEATURE_AND_1_out;
	wire FEATURE_AND_10_out;
	wire FEATURE_AND_2_out;
	wire FEATURE_AND_3_out;
	wire FEATURE_AND_4_out;
	wire FEATURE_AND_5_out;
	wire FEATURE_AND_6_out;
	wire FEATURE_AND_7_out;
	wire FEATURE_AND_8_out;
	wire FEATURE_AND_9_out;
	wire [15:0] MemCore_inst0_output_width_16_num_0;
	wire [15:0] MemCore_inst0_output_width_16_num_1;
	wire [0:0] MemCore_inst0_output_width_1_num_0;
	wire [0:0] MemCore_inst0_output_width_1_num_1;
	wire [0:0] MemCore_inst0_output_width_1_num_2;
	wire [31:0] MemCore_inst0_read_config_data;
	wire [31:0] MemCore_inst0_read_config_data_1;
	wire [7:0] MemCore_inst0_config_1_config_addr_in;
	wire [7:0] MemCore_inst0_config_config_addr_in;
	wire [15:0] SB_ID0_3TRACKS_B16_MemCore_SB_T0_EAST_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_MemCore_SB_T0_NORTH_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_MemCore_SB_T0_SOUTH_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_MemCore_SB_T0_WEST_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_MemCore_SB_T1_EAST_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_MemCore_SB_T1_NORTH_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_MemCore_SB_T1_SOUTH_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_MemCore_SB_T1_WEST_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_MemCore_SB_T2_EAST_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_MemCore_SB_T2_NORTH_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_MemCore_SB_T2_SOUTH_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_MemCore_SB_T2_WEST_SB_OUT_B16;
	wire [31:0] SB_ID0_3TRACKS_B16_MemCore_read_config_data;
	wire [7:0] SB_ID0_3TRACKS_B16_MemCore_config_config_addr_in;
	wire [0:0] SB_ID0_3TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1;
	wire [31:0] SB_ID0_3TRACKS_B1_MemCore_read_config_data;
	wire [7:0] SB_ID0_3TRACKS_B1_MemCore_config_config_addr_in;
	wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T0_EAST_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T0_NORTH_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T0_SOUTH_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T0_WEST_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T1_EAST_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T1_NORTH_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T1_SOUTH_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T1_WEST_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T2_EAST_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T2_NORTH_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T2_SOUTH_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T2_WEST_SB_IN_B16_O;
	wire and_inst0_out;
	wire and_inst1_out;
	wire [7:0] const_0_8_out;
	wire [8:0] const_511_9_out;
	wire coreir_eq_16_inst0_out;
	wire [31:0] read_config_data_or_inst0_out;
	wire [31:0] read_data_mux_O;
	wire [7:0] read_data_mux_S_in;
	wire [31:0] self_config_config_addr_out;
// diodes are put to prevent antenna violations on abutted pins
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T0 (.DIODE(tile_id[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T1 (.DIODE(tile_id[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T2 (.DIODE(tile_id[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T3 (.DIODE(tile_id[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T4 (.DIODE(tile_id[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T5 (.DIODE(tile_id[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T6 (.DIODE(tile_id[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T7 (.DIODE(tile_id[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T8 (.DIODE(tile_id[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T9 (.DIODE(tile_id[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T10 (.DIODE(tile_id[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T11 (.DIODE(tile_id[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T12 (.DIODE(tile_id[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T13 (.DIODE(tile_id[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T14 (.DIODE(tile_id[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T15 (.DIODE(tile_id[15]));
// [start] input diodes
sky130_fd_sc_hd__diode_2 POHAN_DIODE_0 (.DIODE(SB_T0_EAST_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_1 (.DIODE(SB_T0_EAST_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_2 (.DIODE(SB_T0_EAST_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_3 (.DIODE(SB_T0_EAST_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_4 (.DIODE(SB_T0_EAST_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_5 (.DIODE(SB_T0_EAST_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_6 (.DIODE(SB_T0_EAST_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_7 (.DIODE(SB_T0_EAST_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_8 (.DIODE(SB_T0_EAST_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_9 (.DIODE(SB_T0_EAST_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_10 (.DIODE(SB_T0_EAST_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_11 (.DIODE(SB_T0_EAST_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_12 (.DIODE(SB_T0_EAST_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_13 (.DIODE(SB_T0_EAST_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_14 (.DIODE(SB_T0_EAST_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_15 (.DIODE(SB_T0_EAST_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_16 (.DIODE(SB_T0_EAST_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_17 (.DIODE(SB_T0_NORTH_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_18 (.DIODE(SB_T0_NORTH_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_19 (.DIODE(SB_T0_NORTH_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_20 (.DIODE(SB_T0_NORTH_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_21 (.DIODE(SB_T0_NORTH_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_22 (.DIODE(SB_T0_NORTH_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_23 (.DIODE(SB_T0_NORTH_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_24 (.DIODE(SB_T0_NORTH_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_25 (.DIODE(SB_T0_NORTH_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_26 (.DIODE(SB_T0_NORTH_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_27 (.DIODE(SB_T0_NORTH_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_28 (.DIODE(SB_T0_NORTH_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_29 (.DIODE(SB_T0_NORTH_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_30 (.DIODE(SB_T0_NORTH_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_31 (.DIODE(SB_T0_NORTH_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_32 (.DIODE(SB_T0_NORTH_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_33 (.DIODE(SB_T0_NORTH_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_34 (.DIODE(SB_T0_SOUTH_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_35 (.DIODE(SB_T0_SOUTH_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_36 (.DIODE(SB_T0_SOUTH_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_37 (.DIODE(SB_T0_SOUTH_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_38 (.DIODE(SB_T0_SOUTH_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_39 (.DIODE(SB_T0_SOUTH_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_40 (.DIODE(SB_T0_SOUTH_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_41 (.DIODE(SB_T0_SOUTH_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_42 (.DIODE(SB_T0_SOUTH_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_43 (.DIODE(SB_T0_SOUTH_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_44 (.DIODE(SB_T0_SOUTH_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_45 (.DIODE(SB_T0_SOUTH_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_46 (.DIODE(SB_T0_SOUTH_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_47 (.DIODE(SB_T0_SOUTH_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_48 (.DIODE(SB_T0_SOUTH_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_49 (.DIODE(SB_T0_SOUTH_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_50 (.DIODE(SB_T0_SOUTH_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_51 (.DIODE(SB_T0_WEST_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_52 (.DIODE(SB_T0_WEST_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_53 (.DIODE(SB_T0_WEST_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_54 (.DIODE(SB_T0_WEST_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_55 (.DIODE(SB_T0_WEST_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_56 (.DIODE(SB_T0_WEST_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_57 (.DIODE(SB_T0_WEST_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_58 (.DIODE(SB_T0_WEST_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_59 (.DIODE(SB_T0_WEST_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_60 (.DIODE(SB_T0_WEST_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_61 (.DIODE(SB_T0_WEST_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_62 (.DIODE(SB_T0_WEST_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_63 (.DIODE(SB_T0_WEST_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_64 (.DIODE(SB_T0_WEST_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_65 (.DIODE(SB_T0_WEST_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_66 (.DIODE(SB_T0_WEST_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_67 (.DIODE(SB_T0_WEST_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_68 (.DIODE(SB_T1_EAST_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_69 (.DIODE(SB_T1_EAST_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_70 (.DIODE(SB_T1_EAST_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_71 (.DIODE(SB_T1_EAST_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_72 (.DIODE(SB_T1_EAST_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_73 (.DIODE(SB_T1_EAST_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_74 (.DIODE(SB_T1_EAST_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_75 (.DIODE(SB_T1_EAST_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_76 (.DIODE(SB_T1_EAST_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_77 (.DIODE(SB_T1_EAST_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_78 (.DIODE(SB_T1_EAST_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_79 (.DIODE(SB_T1_EAST_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_80 (.DIODE(SB_T1_EAST_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_81 (.DIODE(SB_T1_EAST_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_82 (.DIODE(SB_T1_EAST_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_83 (.DIODE(SB_T1_EAST_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_84 (.DIODE(SB_T1_EAST_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_85 (.DIODE(SB_T1_NORTH_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_86 (.DIODE(SB_T1_NORTH_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_87 (.DIODE(SB_T1_NORTH_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_88 (.DIODE(SB_T1_NORTH_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_89 (.DIODE(SB_T1_NORTH_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_90 (.DIODE(SB_T1_NORTH_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_91 (.DIODE(SB_T1_NORTH_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_92 (.DIODE(SB_T1_NORTH_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_93 (.DIODE(SB_T1_NORTH_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_94 (.DIODE(SB_T1_NORTH_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_95 (.DIODE(SB_T1_NORTH_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_96 (.DIODE(SB_T1_NORTH_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_97 (.DIODE(SB_T1_NORTH_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_98 (.DIODE(SB_T1_NORTH_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_99 (.DIODE(SB_T1_NORTH_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_100 (.DIODE(SB_T1_NORTH_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_101 (.DIODE(SB_T1_NORTH_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_102 (.DIODE(SB_T1_SOUTH_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_103 (.DIODE(SB_T1_SOUTH_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_104 (.DIODE(SB_T1_SOUTH_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_105 (.DIODE(SB_T1_SOUTH_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_106 (.DIODE(SB_T1_SOUTH_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_107 (.DIODE(SB_T1_SOUTH_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_108 (.DIODE(SB_T1_SOUTH_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_109 (.DIODE(SB_T1_SOUTH_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_110 (.DIODE(SB_T1_SOUTH_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_111 (.DIODE(SB_T1_SOUTH_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_112 (.DIODE(SB_T1_SOUTH_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_113 (.DIODE(SB_T1_SOUTH_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_114 (.DIODE(SB_T1_SOUTH_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_115 (.DIODE(SB_T1_SOUTH_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_116 (.DIODE(SB_T1_SOUTH_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_117 (.DIODE(SB_T1_SOUTH_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_118 (.DIODE(SB_T1_SOUTH_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_119 (.DIODE(SB_T1_WEST_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_120 (.DIODE(SB_T1_WEST_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_121 (.DIODE(SB_T1_WEST_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_122 (.DIODE(SB_T1_WEST_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_123 (.DIODE(SB_T1_WEST_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_124 (.DIODE(SB_T1_WEST_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_125 (.DIODE(SB_T1_WEST_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_126 (.DIODE(SB_T1_WEST_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_127 (.DIODE(SB_T1_WEST_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_128 (.DIODE(SB_T1_WEST_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_129 (.DIODE(SB_T1_WEST_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_130 (.DIODE(SB_T1_WEST_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_131 (.DIODE(SB_T1_WEST_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_132 (.DIODE(SB_T1_WEST_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_133 (.DIODE(SB_T1_WEST_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_134 (.DIODE(SB_T1_WEST_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_135 (.DIODE(SB_T1_WEST_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_136 (.DIODE(SB_T2_EAST_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_137 (.DIODE(SB_T2_EAST_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_138 (.DIODE(SB_T2_EAST_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_139 (.DIODE(SB_T2_EAST_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_140 (.DIODE(SB_T2_EAST_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_141 (.DIODE(SB_T2_EAST_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_142 (.DIODE(SB_T2_EAST_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_143 (.DIODE(SB_T2_EAST_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_144 (.DIODE(SB_T2_EAST_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_145 (.DIODE(SB_T2_EAST_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_146 (.DIODE(SB_T2_EAST_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_147 (.DIODE(SB_T2_EAST_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_148 (.DIODE(SB_T2_EAST_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_149 (.DIODE(SB_T2_EAST_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_150 (.DIODE(SB_T2_EAST_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_151 (.DIODE(SB_T2_EAST_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_152 (.DIODE(SB_T2_EAST_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_153 (.DIODE(SB_T2_NORTH_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_154 (.DIODE(SB_T2_NORTH_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_155 (.DIODE(SB_T2_NORTH_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_156 (.DIODE(SB_T2_NORTH_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_157 (.DIODE(SB_T2_NORTH_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_158 (.DIODE(SB_T2_NORTH_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_159 (.DIODE(SB_T2_NORTH_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_160 (.DIODE(SB_T2_NORTH_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_161 (.DIODE(SB_T2_NORTH_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_162 (.DIODE(SB_T2_NORTH_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_163 (.DIODE(SB_T2_NORTH_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_164 (.DIODE(SB_T2_NORTH_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_165 (.DIODE(SB_T2_NORTH_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_166 (.DIODE(SB_T2_NORTH_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_167 (.DIODE(SB_T2_NORTH_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_168 (.DIODE(SB_T2_NORTH_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_169 (.DIODE(SB_T2_NORTH_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_170 (.DIODE(SB_T2_SOUTH_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_171 (.DIODE(SB_T2_SOUTH_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_172 (.DIODE(SB_T2_SOUTH_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_173 (.DIODE(SB_T2_SOUTH_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_174 (.DIODE(SB_T2_SOUTH_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_175 (.DIODE(SB_T2_SOUTH_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_176 (.DIODE(SB_T2_SOUTH_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_177 (.DIODE(SB_T2_SOUTH_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_178 (.DIODE(SB_T2_SOUTH_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_179 (.DIODE(SB_T2_SOUTH_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_180 (.DIODE(SB_T2_SOUTH_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_181 (.DIODE(SB_T2_SOUTH_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_182 (.DIODE(SB_T2_SOUTH_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_183 (.DIODE(SB_T2_SOUTH_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_184 (.DIODE(SB_T2_SOUTH_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_185 (.DIODE(SB_T2_SOUTH_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_186 (.DIODE(SB_T2_SOUTH_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_187 (.DIODE(SB_T2_WEST_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_188 (.DIODE(SB_T2_WEST_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_189 (.DIODE(SB_T2_WEST_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_190 (.DIODE(SB_T2_WEST_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_191 (.DIODE(SB_T2_WEST_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_192 (.DIODE(SB_T2_WEST_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_193 (.DIODE(SB_T2_WEST_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_194 (.DIODE(SB_T2_WEST_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_195 (.DIODE(SB_T2_WEST_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_196 (.DIODE(SB_T2_WEST_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_197 (.DIODE(SB_T2_WEST_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_198 (.DIODE(SB_T2_WEST_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_199 (.DIODE(SB_T2_WEST_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_200 (.DIODE(SB_T2_WEST_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_201 (.DIODE(SB_T2_WEST_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_202 (.DIODE(SB_T2_WEST_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_203 (.DIODE(SB_T2_WEST_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_204 (.DIODE(clk));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_205 (.DIODE(clk_pass_through));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_206 (.DIODE(config_config_addr[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_207 (.DIODE(config_config_addr[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_208 (.DIODE(config_config_addr[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_209 (.DIODE(config_config_addr[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_210 (.DIODE(config_config_addr[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_211 (.DIODE(config_config_addr[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_212 (.DIODE(config_config_addr[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_213 (.DIODE(config_config_addr[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_214 (.DIODE(config_config_addr[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_215 (.DIODE(config_config_addr[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_216 (.DIODE(config_config_addr[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_217 (.DIODE(config_config_addr[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_218 (.DIODE(config_config_addr[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_219 (.DIODE(config_config_addr[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_220 (.DIODE(config_config_addr[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_221 (.DIODE(config_config_addr[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_222 (.DIODE(config_config_addr[16]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_223 (.DIODE(config_config_addr[17]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_224 (.DIODE(config_config_addr[18]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_225 (.DIODE(config_config_addr[19]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_226 (.DIODE(config_config_addr[20]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_227 (.DIODE(config_config_addr[21]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_228 (.DIODE(config_config_addr[22]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_229 (.DIODE(config_config_addr[23]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_230 (.DIODE(config_config_addr[24]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_231 (.DIODE(config_config_addr[25]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_232 (.DIODE(config_config_addr[26]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_233 (.DIODE(config_config_addr[27]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_234 (.DIODE(config_config_addr[28]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_235 (.DIODE(config_config_addr[29]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_236 (.DIODE(config_config_addr[30]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_237 (.DIODE(config_config_addr[31]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_238 (.DIODE(config_config_data[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_239 (.DIODE(config_config_data[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_240 (.DIODE(config_config_data[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_241 (.DIODE(config_config_data[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_242 (.DIODE(config_config_data[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_243 (.DIODE(config_config_data[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_244 (.DIODE(config_config_data[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_245 (.DIODE(config_config_data[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_246 (.DIODE(config_config_data[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_247 (.DIODE(config_config_data[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_248 (.DIODE(config_config_data[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_249 (.DIODE(config_config_data[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_250 (.DIODE(config_config_data[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_251 (.DIODE(config_config_data[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_252 (.DIODE(config_config_data[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_253 (.DIODE(config_config_data[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_254 (.DIODE(config_config_data[16]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_255 (.DIODE(config_config_data[17]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_256 (.DIODE(config_config_data[18]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_257 (.DIODE(config_config_data[19]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_258 (.DIODE(config_config_data[20]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_259 (.DIODE(config_config_data[21]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_260 (.DIODE(config_config_data[22]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_261 (.DIODE(config_config_data[23]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_262 (.DIODE(config_config_data[24]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_263 (.DIODE(config_config_data[25]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_264 (.DIODE(config_config_data[26]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_265 (.DIODE(config_config_data[27]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_266 (.DIODE(config_config_data[28]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_267 (.DIODE(config_config_data[29]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_268 (.DIODE(config_config_data[30]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_269 (.DIODE(config_config_data[31]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_270 (.DIODE(config_read[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_271 (.DIODE(config_write[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_272 (.DIODE(read_config_data_in[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_273 (.DIODE(read_config_data_in[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_274 (.DIODE(read_config_data_in[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_275 (.DIODE(read_config_data_in[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_276 (.DIODE(read_config_data_in[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_277 (.DIODE(read_config_data_in[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_278 (.DIODE(read_config_data_in[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_279 (.DIODE(read_config_data_in[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_280 (.DIODE(read_config_data_in[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_281 (.DIODE(read_config_data_in[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_282 (.DIODE(read_config_data_in[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_283 (.DIODE(read_config_data_in[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_284 (.DIODE(read_config_data_in[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_285 (.DIODE(read_config_data_in[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_286 (.DIODE(read_config_data_in[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_287 (.DIODE(read_config_data_in[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_288 (.DIODE(read_config_data_in[16]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_289 (.DIODE(read_config_data_in[17]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_290 (.DIODE(read_config_data_in[18]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_291 (.DIODE(read_config_data_in[19]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_292 (.DIODE(read_config_data_in[20]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_293 (.DIODE(read_config_data_in[21]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_294 (.DIODE(read_config_data_in[22]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_295 (.DIODE(read_config_data_in[23]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_296 (.DIODE(read_config_data_in[24]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_297 (.DIODE(read_config_data_in[25]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_298 (.DIODE(read_config_data_in[26]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_299 (.DIODE(read_config_data_in[27]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_300 (.DIODE(read_config_data_in[28]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_301 (.DIODE(read_config_data_in[29]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_302 (.DIODE(read_config_data_in[30]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_303 (.DIODE(read_config_data_in[31]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_304 (.DIODE(reset));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_305 (.DIODE(stall[0]));
// [end] input diodes

// [start] output diodes
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_306 (.DIODE(SB_T0_EAST_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_307 (.DIODE(SB_T0_EAST_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_308 (.DIODE(SB_T0_EAST_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_309 (.DIODE(SB_T0_EAST_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_310 (.DIODE(SB_T0_EAST_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_311 (.DIODE(SB_T0_EAST_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_312 (.DIODE(SB_T0_EAST_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_313 (.DIODE(SB_T0_EAST_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_314 (.DIODE(SB_T0_EAST_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_315 (.DIODE(SB_T0_EAST_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_316 (.DIODE(SB_T0_EAST_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_317 (.DIODE(SB_T0_EAST_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_318 (.DIODE(SB_T0_EAST_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_319 (.DIODE(SB_T0_EAST_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_320 (.DIODE(SB_T0_EAST_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_321 (.DIODE(SB_T0_EAST_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_322 (.DIODE(SB_T0_EAST_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_323 (.DIODE(SB_T0_NORTH_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_324 (.DIODE(SB_T0_NORTH_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_325 (.DIODE(SB_T0_NORTH_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_326 (.DIODE(SB_T0_NORTH_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_327 (.DIODE(SB_T0_NORTH_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_328 (.DIODE(SB_T0_NORTH_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_329 (.DIODE(SB_T0_NORTH_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_330 (.DIODE(SB_T0_NORTH_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_331 (.DIODE(SB_T0_NORTH_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_332 (.DIODE(SB_T0_NORTH_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_333 (.DIODE(SB_T0_NORTH_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_334 (.DIODE(SB_T0_NORTH_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_335 (.DIODE(SB_T0_NORTH_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_336 (.DIODE(SB_T0_NORTH_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_337 (.DIODE(SB_T0_NORTH_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_338 (.DIODE(SB_T0_NORTH_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_339 (.DIODE(SB_T0_NORTH_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_340 (.DIODE(SB_T0_SOUTH_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_341 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_342 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_343 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_344 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_345 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_346 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_347 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_348 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_349 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_350 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_351 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_352 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_353 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_354 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_355 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_356 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_357 (.DIODE(SB_T0_WEST_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_358 (.DIODE(SB_T0_WEST_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_359 (.DIODE(SB_T0_WEST_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_360 (.DIODE(SB_T0_WEST_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_361 (.DIODE(SB_T0_WEST_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_362 (.DIODE(SB_T0_WEST_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_363 (.DIODE(SB_T0_WEST_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_364 (.DIODE(SB_T0_WEST_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_365 (.DIODE(SB_T0_WEST_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_366 (.DIODE(SB_T0_WEST_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_367 (.DIODE(SB_T0_WEST_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_368 (.DIODE(SB_T0_WEST_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_369 (.DIODE(SB_T0_WEST_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_370 (.DIODE(SB_T0_WEST_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_371 (.DIODE(SB_T0_WEST_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_372 (.DIODE(SB_T0_WEST_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_373 (.DIODE(SB_T0_WEST_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_374 (.DIODE(SB_T1_EAST_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_375 (.DIODE(SB_T1_EAST_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_376 (.DIODE(SB_T1_EAST_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_377 (.DIODE(SB_T1_EAST_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_378 (.DIODE(SB_T1_EAST_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_379 (.DIODE(SB_T1_EAST_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_380 (.DIODE(SB_T1_EAST_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_381 (.DIODE(SB_T1_EAST_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_382 (.DIODE(SB_T1_EAST_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_383 (.DIODE(SB_T1_EAST_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_384 (.DIODE(SB_T1_EAST_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_385 (.DIODE(SB_T1_EAST_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_386 (.DIODE(SB_T1_EAST_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_387 (.DIODE(SB_T1_EAST_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_388 (.DIODE(SB_T1_EAST_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_389 (.DIODE(SB_T1_EAST_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_390 (.DIODE(SB_T1_EAST_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_391 (.DIODE(SB_T1_NORTH_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_392 (.DIODE(SB_T1_NORTH_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_393 (.DIODE(SB_T1_NORTH_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_394 (.DIODE(SB_T1_NORTH_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_395 (.DIODE(SB_T1_NORTH_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_396 (.DIODE(SB_T1_NORTH_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_397 (.DIODE(SB_T1_NORTH_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_398 (.DIODE(SB_T1_NORTH_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_399 (.DIODE(SB_T1_NORTH_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_400 (.DIODE(SB_T1_NORTH_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_401 (.DIODE(SB_T1_NORTH_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_402 (.DIODE(SB_T1_NORTH_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_403 (.DIODE(SB_T1_NORTH_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_404 (.DIODE(SB_T1_NORTH_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_405 (.DIODE(SB_T1_NORTH_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_406 (.DIODE(SB_T1_NORTH_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_407 (.DIODE(SB_T1_NORTH_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_408 (.DIODE(SB_T1_SOUTH_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_409 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_410 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_411 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_412 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_413 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_414 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_415 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_416 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_417 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_418 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_419 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_420 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_421 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_422 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_423 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_424 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_425 (.DIODE(SB_T1_WEST_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_426 (.DIODE(SB_T1_WEST_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_427 (.DIODE(SB_T1_WEST_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_428 (.DIODE(SB_T1_WEST_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_429 (.DIODE(SB_T1_WEST_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_430 (.DIODE(SB_T1_WEST_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_431 (.DIODE(SB_T1_WEST_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_432 (.DIODE(SB_T1_WEST_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_433 (.DIODE(SB_T1_WEST_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_434 (.DIODE(SB_T1_WEST_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_435 (.DIODE(SB_T1_WEST_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_436 (.DIODE(SB_T1_WEST_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_437 (.DIODE(SB_T1_WEST_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_438 (.DIODE(SB_T1_WEST_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_439 (.DIODE(SB_T1_WEST_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_440 (.DIODE(SB_T1_WEST_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_441 (.DIODE(SB_T1_WEST_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_442 (.DIODE(SB_T2_EAST_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_443 (.DIODE(SB_T2_EAST_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_444 (.DIODE(SB_T2_EAST_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_445 (.DIODE(SB_T2_EAST_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_446 (.DIODE(SB_T2_EAST_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_447 (.DIODE(SB_T2_EAST_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_448 (.DIODE(SB_T2_EAST_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_449 (.DIODE(SB_T2_EAST_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_450 (.DIODE(SB_T2_EAST_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_451 (.DIODE(SB_T2_EAST_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_452 (.DIODE(SB_T2_EAST_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_453 (.DIODE(SB_T2_EAST_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_454 (.DIODE(SB_T2_EAST_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_455 (.DIODE(SB_T2_EAST_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_456 (.DIODE(SB_T2_EAST_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_457 (.DIODE(SB_T2_EAST_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_458 (.DIODE(SB_T2_EAST_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_459 (.DIODE(SB_T2_NORTH_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_460 (.DIODE(SB_T2_NORTH_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_461 (.DIODE(SB_T2_NORTH_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_462 (.DIODE(SB_T2_NORTH_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_463 (.DIODE(SB_T2_NORTH_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_464 (.DIODE(SB_T2_NORTH_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_465 (.DIODE(SB_T2_NORTH_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_466 (.DIODE(SB_T2_NORTH_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_467 (.DIODE(SB_T2_NORTH_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_468 (.DIODE(SB_T2_NORTH_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_469 (.DIODE(SB_T2_NORTH_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_470 (.DIODE(SB_T2_NORTH_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_471 (.DIODE(SB_T2_NORTH_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_472 (.DIODE(SB_T2_NORTH_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_473 (.DIODE(SB_T2_NORTH_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_474 (.DIODE(SB_T2_NORTH_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_475 (.DIODE(SB_T2_NORTH_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_476 (.DIODE(SB_T2_SOUTH_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_477 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_478 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_479 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_480 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_481 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_482 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_483 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_484 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_485 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_486 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_487 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_488 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_489 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_490 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_491 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_492 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_493 (.DIODE(SB_T2_WEST_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_494 (.DIODE(SB_T2_WEST_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_495 (.DIODE(SB_T2_WEST_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_496 (.DIODE(SB_T2_WEST_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_497 (.DIODE(SB_T2_WEST_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_498 (.DIODE(SB_T2_WEST_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_499 (.DIODE(SB_T2_WEST_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_500 (.DIODE(SB_T2_WEST_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_501 (.DIODE(SB_T2_WEST_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_502 (.DIODE(SB_T2_WEST_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_503 (.DIODE(SB_T2_WEST_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_504 (.DIODE(SB_T2_WEST_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_505 (.DIODE(SB_T2_WEST_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_506 (.DIODE(SB_T2_WEST_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_507 (.DIODE(SB_T2_WEST_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_508 (.DIODE(SB_T2_WEST_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_509 (.DIODE(SB_T2_WEST_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_510 (.DIODE(clk_out));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_511 (.DIODE(clk_pass_through_out_bot));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_512 (.DIODE(config_out_config_addr[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_513 (.DIODE(config_out_config_addr[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_514 (.DIODE(config_out_config_addr[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_515 (.DIODE(config_out_config_addr[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_516 (.DIODE(config_out_config_addr[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_517 (.DIODE(config_out_config_addr[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_518 (.DIODE(config_out_config_addr[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_519 (.DIODE(config_out_config_addr[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_520 (.DIODE(config_out_config_addr[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_521 (.DIODE(config_out_config_addr[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_522 (.DIODE(config_out_config_addr[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_523 (.DIODE(config_out_config_addr[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_524 (.DIODE(config_out_config_addr[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_525 (.DIODE(config_out_config_addr[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_526 (.DIODE(config_out_config_addr[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_527 (.DIODE(config_out_config_addr[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_528 (.DIODE(config_out_config_addr[16]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_529 (.DIODE(config_out_config_addr[17]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_530 (.DIODE(config_out_config_addr[18]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_531 (.DIODE(config_out_config_addr[19]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_532 (.DIODE(config_out_config_addr[20]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_533 (.DIODE(config_out_config_addr[21]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_534 (.DIODE(config_out_config_addr[22]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_535 (.DIODE(config_out_config_addr[23]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_536 (.DIODE(config_out_config_addr[24]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_537 (.DIODE(config_out_config_addr[25]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_538 (.DIODE(config_out_config_addr[26]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_539 (.DIODE(config_out_config_addr[27]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_540 (.DIODE(config_out_config_addr[28]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_541 (.DIODE(config_out_config_addr[29]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_542 (.DIODE(config_out_config_addr[30]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_543 (.DIODE(config_out_config_addr[31]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_544 (.DIODE(config_out_config_data[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_545 (.DIODE(config_out_config_data[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_546 (.DIODE(config_out_config_data[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_547 (.DIODE(config_out_config_data[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_548 (.DIODE(config_out_config_data[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_549 (.DIODE(config_out_config_data[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_550 (.DIODE(config_out_config_data[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_551 (.DIODE(config_out_config_data[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_552 (.DIODE(config_out_config_data[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_553 (.DIODE(config_out_config_data[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_554 (.DIODE(config_out_config_data[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_555 (.DIODE(config_out_config_data[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_556 (.DIODE(config_out_config_data[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_557 (.DIODE(config_out_config_data[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_558 (.DIODE(config_out_config_data[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_559 (.DIODE(config_out_config_data[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_560 (.DIODE(config_out_config_data[16]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_561 (.DIODE(config_out_config_data[17]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_562 (.DIODE(config_out_config_data[18]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_563 (.DIODE(config_out_config_data[19]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_564 (.DIODE(config_out_config_data[20]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_565 (.DIODE(config_out_config_data[21]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_566 (.DIODE(config_out_config_data[22]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_567 (.DIODE(config_out_config_data[23]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_568 (.DIODE(config_out_config_data[24]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_569 (.DIODE(config_out_config_data[25]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_570 (.DIODE(config_out_config_data[26]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_571 (.DIODE(config_out_config_data[27]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_572 (.DIODE(config_out_config_data[28]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_573 (.DIODE(config_out_config_data[29]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_574 (.DIODE(config_out_config_data[30]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_575 (.DIODE(config_out_config_data[31]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_576 (.DIODE(config_out_read[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_577 (.DIODE(config_out_write[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_578 (.DIODE(read_config_data[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_579 (.DIODE(read_config_data[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_580 (.DIODE(read_config_data[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_581 (.DIODE(read_config_data[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_582 (.DIODE(read_config_data[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_583 (.DIODE(read_config_data[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_584 (.DIODE(read_config_data[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_585 (.DIODE(read_config_data[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_586 (.DIODE(read_config_data[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_587 (.DIODE(read_config_data[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_588 (.DIODE(read_config_data[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_589 (.DIODE(read_config_data[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_590 (.DIODE(read_config_data[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_591 (.DIODE(read_config_data[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_592 (.DIODE(read_config_data[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_593 (.DIODE(read_config_data[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_594 (.DIODE(read_config_data[16]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_595 (.DIODE(read_config_data[17]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_596 (.DIODE(read_config_data[18]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_597 (.DIODE(read_config_data[19]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_598 (.DIODE(read_config_data[20]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_599 (.DIODE(read_config_data[21]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_600 (.DIODE(read_config_data[22]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_601 (.DIODE(read_config_data[23]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_602 (.DIODE(read_config_data[24]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_603 (.DIODE(read_config_data[25]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_604 (.DIODE(read_config_data[26]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_605 (.DIODE(read_config_data[27]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_606 (.DIODE(read_config_data[28]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_607 (.DIODE(read_config_data[29]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_608 (.DIODE(read_config_data[30]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_609 (.DIODE(read_config_data[31]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_610 (.DIODE(reset_out));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_611 (.DIODE(stall_out[0]));
// [end] output diodes
	CB_flush CB_flush(
		.I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
		.I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
		.I_10(WIRE_SB_T2_EAST_SB_IN_B1_O),
		.I_11(WIRE_SB_T2_WEST_SB_IN_B1_O),
		.I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
		.I_3(WIRE_SB_T0_WEST_SB_IN_B1_O),
		.I_4(WIRE_SB_T1_NORTH_SB_IN_B1_O),
		.I_5(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
		.I_6(WIRE_SB_T1_EAST_SB_IN_B1_O),
		.I_7(WIRE_SB_T1_WEST_SB_IN_B1_O),
		.I_8(WIRE_SB_T2_NORTH_SB_IN_B1_O),
		.I_9(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
		.O(CB_flush_O),
		.clk(clk),
		.config_config_addr(CB_flush_config_config_addr_in),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_2_out),
		.read_config_data(CB_flush_read_config_data),
		.reset(reset)
	);
	mantle_wire__typeBitIn8 CB_flush_config_config_addr(
		.in(CB_flush_config_config_addr_in),
		.out(self_config_config_addr_out[31:24])
	);
	CB_input_width_16_num_0 CB_input_width_16_num_0(
		.I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
		.I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
		.I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
		.I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
		.I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
		.I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
		.I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
		.I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
		.I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
		.I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
		.I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
		.I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
		.O(CB_input_width_16_num_0_O),
		.clk(clk),
		.config_config_addr(CB_input_width_16_num_0_config_config_addr_in),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_3_out),
		.read_config_data(CB_input_width_16_num_0_read_config_data),
		.reset(reset)
	);
	mantle_wire__typeBitIn8 CB_input_width_16_num_0_config_config_addr(
		.in(CB_input_width_16_num_0_config_config_addr_in),
		.out(self_config_config_addr_out[31:24])
	);
	CB_input_width_16_num_1 CB_input_width_16_num_1(
		.I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
		.I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
		.I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
		.I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
		.I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
		.I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
		.I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
		.I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
		.I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
		.I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
		.I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
		.I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
		.O(CB_input_width_16_num_1_O),
		.clk(clk),
		.config_config_addr(CB_input_width_16_num_1_config_config_addr_in),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_4_out),
		.read_config_data(CB_input_width_16_num_1_read_config_data),
		.reset(reset)
	);
	mantle_wire__typeBitIn8 CB_input_width_16_num_1_config_config_addr(
		.in(CB_input_width_16_num_1_config_config_addr_in),
		.out(self_config_config_addr_out[31:24])
	);
	CB_input_width_16_num_2 CB_input_width_16_num_2(
		.I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
		.I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
		.I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
		.I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
		.I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
		.I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
		.I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
		.I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
		.I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
		.I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
		.I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
		.I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
		.O(CB_input_width_16_num_2_O),
		.clk(clk),
		.config_config_addr(CB_input_width_16_num_2_config_config_addr_in),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_5_out),
		.read_config_data(CB_input_width_16_num_2_read_config_data),
		.reset(reset)
	);
	mantle_wire__typeBitIn8 CB_input_width_16_num_2_config_config_addr(
		.in(CB_input_width_16_num_2_config_config_addr_in),
		.out(self_config_config_addr_out[31:24])
	);
	CB_input_width_16_num_3 CB_input_width_16_num_3(
		.I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
		.I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
		.I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
		.I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
		.I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
		.I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
		.I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
		.I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
		.I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
		.I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
		.I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
		.I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
		.O(CB_input_width_16_num_3_O),
		.clk(clk),
		.config_config_addr(CB_input_width_16_num_3_config_config_addr_in),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_6_out),
		.read_config_data(CB_input_width_16_num_3_read_config_data),
		.reset(reset)
	);
	mantle_wire__typeBitIn8 CB_input_width_16_num_3_config_config_addr(
		.in(CB_input_width_16_num_3_config_config_addr_in),
		.out(self_config_config_addr_out[31:24])
	);
	CB_input_width_1_num_0 CB_input_width_1_num_0(
		.I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
		.I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
		.I_10(WIRE_SB_T2_EAST_SB_IN_B1_O),
		.I_11(WIRE_SB_T2_WEST_SB_IN_B1_O),
		.I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
		.I_3(WIRE_SB_T0_WEST_SB_IN_B1_O),
		.I_4(WIRE_SB_T1_NORTH_SB_IN_B1_O),
		.I_5(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
		.I_6(WIRE_SB_T1_EAST_SB_IN_B1_O),
		.I_7(WIRE_SB_T1_WEST_SB_IN_B1_O),
		.I_8(WIRE_SB_T2_NORTH_SB_IN_B1_O),
		.I_9(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
		.O(CB_input_width_1_num_0_O),
		.clk(clk),
		.config_config_addr(CB_input_width_1_num_0_config_config_addr_in),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_7_out),
		.read_config_data(CB_input_width_1_num_0_read_config_data),
		.reset(reset)
	);
	mantle_wire__typeBitIn8 CB_input_width_1_num_0_config_config_addr(
		.in(CB_input_width_1_num_0_config_config_addr_in),
		.out(self_config_config_addr_out[31:24])
	);
	CB_input_width_1_num_1 CB_input_width_1_num_1(
		.I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
		.I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
		.I_10(WIRE_SB_T2_EAST_SB_IN_B1_O),
		.I_11(WIRE_SB_T2_WEST_SB_IN_B1_O),
		.I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
		.I_3(WIRE_SB_T0_WEST_SB_IN_B1_O),
		.I_4(WIRE_SB_T1_NORTH_SB_IN_B1_O),
		.I_5(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
		.I_6(WIRE_SB_T1_EAST_SB_IN_B1_O),
		.I_7(WIRE_SB_T1_WEST_SB_IN_B1_O),
		.I_8(WIRE_SB_T2_NORTH_SB_IN_B1_O),
		.I_9(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
		.O(CB_input_width_1_num_1_O),
		.clk(clk),
		.config_config_addr(CB_input_width_1_num_1_config_config_addr_in),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_8_out),
		.read_config_data(CB_input_width_1_num_1_read_config_data),
		.reset(reset)
	);
	mantle_wire__typeBitIn8 CB_input_width_1_num_1_config_config_addr(
		.in(CB_input_width_1_num_1_config_config_addr_in),
		.out(self_config_config_addr_out[31:24])
	);
	Decode08 DECODE_FEATURE_0(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_0_O)
	);
	Decode18 DECODE_FEATURE_1(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_1_O)
	);
	Decode108 DECODE_FEATURE_10(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_10_O)
	);
	Decode28 DECODE_FEATURE_2(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_2_O)
	);
	Decode38 DECODE_FEATURE_3(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_3_O)
	);
	Decode48 DECODE_FEATURE_4(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_4_O)
	);
	Decode58 DECODE_FEATURE_5(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_5_O)
	);
	Decode68 DECODE_FEATURE_6(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_6_O)
	);
	Decode78 DECODE_FEATURE_7(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_7_O)
	);
	Decode88 DECODE_FEATURE_8(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_8_O)
	);
	Decode98 DECODE_FEATURE_9(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_9_O)
	);
	corebit_and FEATURE_AND_0(
		.in0(DECODE_FEATURE_0_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_0_out)
	);
	corebit_and FEATURE_AND_1(
		.in0(DECODE_FEATURE_1_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_1_out)
	);
	corebit_and FEATURE_AND_10(
		.in0(DECODE_FEATURE_10_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_10_out)
	);
	corebit_and FEATURE_AND_2(
		.in0(DECODE_FEATURE_2_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_2_out)
	);
	corebit_and FEATURE_AND_3(
		.in0(DECODE_FEATURE_3_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_3_out)
	);
	corebit_and FEATURE_AND_4(
		.in0(DECODE_FEATURE_4_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_4_out)
	);
	corebit_and FEATURE_AND_5(
		.in0(DECODE_FEATURE_5_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_5_out)
	);
	corebit_and FEATURE_AND_6(
		.in0(DECODE_FEATURE_6_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_6_out)
	);
	corebit_and FEATURE_AND_7(
		.in0(DECODE_FEATURE_7_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_7_out)
	);
	corebit_and FEATURE_AND_8(
		.in0(DECODE_FEATURE_8_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_8_out)
	);
	corebit_and FEATURE_AND_9(
		.in0(DECODE_FEATURE_9_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_9_out)
	);
	MemCore MemCore_inst0(
		.clk(clk),
		.config_1_config_addr(MemCore_inst0_config_1_config_addr_in),
		.config_1_config_data(config_config_data),
		.config_1_read(config_read),
		.config_1_write(FEATURE_AND_1_out),
		.config_config_addr(MemCore_inst0_config_config_addr_in),
		.config_config_data(config_config_data),
		.config_en_0(DECODE_FEATURE_1_O),
		.config_read(config_read),
		.config_write(FEATURE_AND_0_out),
		.flush(CB_flush_O),
		.input_width_16_num_0(CB_input_width_16_num_0_O),
		.input_width_16_num_1(CB_input_width_16_num_1_O),
		.input_width_16_num_2(CB_input_width_16_num_2_O),
		.input_width_16_num_3(CB_input_width_16_num_3_O),
		.input_width_1_num_0(CB_input_width_1_num_0_O),
		.input_width_1_num_1(CB_input_width_1_num_1_O),
		.output_width_16_num_0(MemCore_inst0_output_width_16_num_0),
		.output_width_16_num_1(MemCore_inst0_output_width_16_num_1),
		.output_width_1_num_0(MemCore_inst0_output_width_1_num_0),
		.output_width_1_num_1(MemCore_inst0_output_width_1_num_1),
		.output_width_1_num_2(MemCore_inst0_output_width_1_num_2),
		.read_config_data(MemCore_inst0_read_config_data),
		.read_config_data_1(MemCore_inst0_read_config_data_1),
		.reset(reset),
		.stall(stall)
	);
	mantle_wire__typeBitIn8 MemCore_inst0_config_1_config_addr(
		.in(MemCore_inst0_config_1_config_addr_in),
		.out(self_config_config_addr_out[31:24])
	);
	mantle_wire__typeBitIn8 MemCore_inst0_config_config_addr(
		.in(MemCore_inst0_config_config_addr_in),
		.out(self_config_config_addr_out[31:24])
	);
	SB_ID0_3TRACKS_B16_MemCore SB_ID0_3TRACKS_B16_MemCore(
		.SB_T0_EAST_SB_IN_B16(SB_T0_EAST_SB_IN_B16),
		.SB_T0_EAST_SB_OUT_B16(SB_ID0_3TRACKS_B16_MemCore_SB_T0_EAST_SB_OUT_B16),
		.SB_T0_NORTH_SB_IN_B16(SB_T0_NORTH_SB_IN_B16),
		.SB_T0_NORTH_SB_OUT_B16(SB_ID0_3TRACKS_B16_MemCore_SB_T0_NORTH_SB_OUT_B16),
		.SB_T0_SOUTH_SB_IN_B16(SB_T0_SOUTH_SB_IN_B16),
		.SB_T0_SOUTH_SB_OUT_B16(SB_ID0_3TRACKS_B16_MemCore_SB_T0_SOUTH_SB_OUT_B16),
		.SB_T0_WEST_SB_IN_B16(SB_T0_WEST_SB_IN_B16),
		.SB_T0_WEST_SB_OUT_B16(SB_ID0_3TRACKS_B16_MemCore_SB_T0_WEST_SB_OUT_B16),
		.SB_T1_EAST_SB_IN_B16(SB_T1_EAST_SB_IN_B16),
		.SB_T1_EAST_SB_OUT_B16(SB_ID0_3TRACKS_B16_MemCore_SB_T1_EAST_SB_OUT_B16),
		.SB_T1_NORTH_SB_IN_B16(SB_T1_NORTH_SB_IN_B16),
		.SB_T1_NORTH_SB_OUT_B16(SB_ID0_3TRACKS_B16_MemCore_SB_T1_NORTH_SB_OUT_B16),
		.SB_T1_SOUTH_SB_IN_B16(SB_T1_SOUTH_SB_IN_B16),
		.SB_T1_SOUTH_SB_OUT_B16(SB_ID0_3TRACKS_B16_MemCore_SB_T1_SOUTH_SB_OUT_B16),
		.SB_T1_WEST_SB_IN_B16(SB_T1_WEST_SB_IN_B16),
		.SB_T1_WEST_SB_OUT_B16(SB_ID0_3TRACKS_B16_MemCore_SB_T1_WEST_SB_OUT_B16),
		.SB_T2_EAST_SB_IN_B16(SB_T2_EAST_SB_IN_B16),
		.SB_T2_EAST_SB_OUT_B16(SB_ID0_3TRACKS_B16_MemCore_SB_T2_EAST_SB_OUT_B16),
		.SB_T2_NORTH_SB_IN_B16(SB_T2_NORTH_SB_IN_B16),
		.SB_T2_NORTH_SB_OUT_B16(SB_ID0_3TRACKS_B16_MemCore_SB_T2_NORTH_SB_OUT_B16),
		.SB_T2_SOUTH_SB_IN_B16(SB_T2_SOUTH_SB_IN_B16),
		.SB_T2_SOUTH_SB_OUT_B16(SB_ID0_3TRACKS_B16_MemCore_SB_T2_SOUTH_SB_OUT_B16),
		.SB_T2_WEST_SB_IN_B16(SB_T2_WEST_SB_IN_B16),
		.SB_T2_WEST_SB_OUT_B16(SB_ID0_3TRACKS_B16_MemCore_SB_T2_WEST_SB_OUT_B16),
		.clk(clk),
		.config_config_addr(SB_ID0_3TRACKS_B16_MemCore_config_config_addr_in),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_10_out),
		.output_width_16_num_0(MemCore_inst0_output_width_16_num_0),
		.output_width_16_num_1(MemCore_inst0_output_width_16_num_1),
		.read_config_data(SB_ID0_3TRACKS_B16_MemCore_read_config_data),
		.reset(reset),
		.stall(stall)
	);
	mantle_wire__typeBitIn8 SB_ID0_3TRACKS_B16_MemCore_config_config_addr(
		.in(SB_ID0_3TRACKS_B16_MemCore_config_config_addr_in),
		.out(self_config_config_addr_out[31:24])
	);
	SB_ID0_3TRACKS_B1_MemCore SB_ID0_3TRACKS_B1_MemCore(
		.SB_T0_EAST_SB_IN_B1(SB_T0_EAST_SB_IN_B1),
		.SB_T0_EAST_SB_OUT_B1(SB_ID0_3TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_NORTH_SB_IN_B1(SB_T0_NORTH_SB_IN_B1),
		.SB_T0_NORTH_SB_OUT_B1(SB_ID0_3TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_IN_B1(SB_T0_SOUTH_SB_IN_B1),
		.SB_T0_SOUTH_SB_OUT_B1(SB_ID0_3TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_WEST_SB_IN_B1(SB_T0_WEST_SB_IN_B1),
		.SB_T0_WEST_SB_OUT_B1(SB_ID0_3TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1),
		.SB_T1_EAST_SB_IN_B1(SB_T1_EAST_SB_IN_B1),
		.SB_T1_EAST_SB_OUT_B1(SB_ID0_3TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_NORTH_SB_IN_B1(SB_T1_NORTH_SB_IN_B1),
		.SB_T1_NORTH_SB_OUT_B1(SB_ID0_3TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_IN_B1(SB_T1_SOUTH_SB_IN_B1),
		.SB_T1_SOUTH_SB_OUT_B1(SB_ID0_3TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_WEST_SB_IN_B1(SB_T1_WEST_SB_IN_B1),
		.SB_T1_WEST_SB_OUT_B1(SB_ID0_3TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1),
		.SB_T2_EAST_SB_IN_B1(SB_T2_EAST_SB_IN_B1),
		.SB_T2_EAST_SB_OUT_B1(SB_ID0_3TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_NORTH_SB_IN_B1(SB_T2_NORTH_SB_IN_B1),
		.SB_T2_NORTH_SB_OUT_B1(SB_ID0_3TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_IN_B1(SB_T2_SOUTH_SB_IN_B1),
		.SB_T2_SOUTH_SB_OUT_B1(SB_ID0_3TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_WEST_SB_IN_B1(SB_T2_WEST_SB_IN_B1),
		.SB_T2_WEST_SB_OUT_B1(SB_ID0_3TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1),
		.clk(clk),
		.config_config_addr(SB_ID0_3TRACKS_B1_MemCore_config_config_addr_in),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_9_out),
		.output_width_1_num_0(MemCore_inst0_output_width_1_num_0),
		.output_width_1_num_1(MemCore_inst0_output_width_1_num_1),
		.output_width_1_num_2(MemCore_inst0_output_width_1_num_2),
		.read_config_data(SB_ID0_3TRACKS_B1_MemCore_read_config_data),
		.reset(reset),
		.stall(stall)
	);
	mantle_wire__typeBitIn8 SB_ID0_3TRACKS_B1_MemCore_config_config_addr(
		.in(SB_ID0_3TRACKS_B1_MemCore_config_config_addr_in),
		.out(self_config_config_addr_out[31:24])
	);
	MuxWrapper_1_1 WIRE_SB_T0_EAST_SB_IN_B1(
		.I(SB_T0_EAST_SB_IN_B1),
		.O(WIRE_SB_T0_EAST_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T0_EAST_SB_IN_B16(
		.I(SB_T0_EAST_SB_IN_B16),
		.O(WIRE_SB_T0_EAST_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T0_NORTH_SB_IN_B1(
		.I(SB_T0_NORTH_SB_IN_B1),
		.O(WIRE_SB_T0_NORTH_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T0_NORTH_SB_IN_B16(
		.I(SB_T0_NORTH_SB_IN_B16),
		.O(WIRE_SB_T0_NORTH_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T0_SOUTH_SB_IN_B1(
		.I(SB_T0_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T0_SOUTH_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T0_SOUTH_SB_IN_B16(
		.I(SB_T0_SOUTH_SB_IN_B16),
		.O(WIRE_SB_T0_SOUTH_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T0_WEST_SB_IN_B1(
		.I(SB_T0_WEST_SB_IN_B1),
		.O(WIRE_SB_T0_WEST_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T0_WEST_SB_IN_B16(
		.I(SB_T0_WEST_SB_IN_B16),
		.O(WIRE_SB_T0_WEST_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T1_EAST_SB_IN_B1(
		.I(SB_T1_EAST_SB_IN_B1),
		.O(WIRE_SB_T1_EAST_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T1_EAST_SB_IN_B16(
		.I(SB_T1_EAST_SB_IN_B16),
		.O(WIRE_SB_T1_EAST_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T1_NORTH_SB_IN_B1(
		.I(SB_T1_NORTH_SB_IN_B1),
		.O(WIRE_SB_T1_NORTH_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T1_NORTH_SB_IN_B16(
		.I(SB_T1_NORTH_SB_IN_B16),
		.O(WIRE_SB_T1_NORTH_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T1_SOUTH_SB_IN_B1(
		.I(SB_T1_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T1_SOUTH_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T1_SOUTH_SB_IN_B16(
		.I(SB_T1_SOUTH_SB_IN_B16),
		.O(WIRE_SB_T1_SOUTH_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T1_WEST_SB_IN_B1(
		.I(SB_T1_WEST_SB_IN_B1),
		.O(WIRE_SB_T1_WEST_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T1_WEST_SB_IN_B16(
		.I(SB_T1_WEST_SB_IN_B16),
		.O(WIRE_SB_T1_WEST_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T2_EAST_SB_IN_B1(
		.I(SB_T2_EAST_SB_IN_B1),
		.O(WIRE_SB_T2_EAST_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T2_EAST_SB_IN_B16(
		.I(SB_T2_EAST_SB_IN_B16),
		.O(WIRE_SB_T2_EAST_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T2_NORTH_SB_IN_B1(
		.I(SB_T2_NORTH_SB_IN_B1),
		.O(WIRE_SB_T2_NORTH_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T2_NORTH_SB_IN_B16(
		.I(SB_T2_NORTH_SB_IN_B16),
		.O(WIRE_SB_T2_NORTH_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T2_SOUTH_SB_IN_B1(
		.I(SB_T2_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T2_SOUTH_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T2_SOUTH_SB_IN_B16(
		.I(SB_T2_SOUTH_SB_IN_B16),
		.O(WIRE_SB_T2_SOUTH_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T2_WEST_SB_IN_B1(
		.I(SB_T2_WEST_SB_IN_B1),
		.O(WIRE_SB_T2_WEST_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T2_WEST_SB_IN_B16(
		.I(SB_T2_WEST_SB_IN_B16),
		.O(WIRE_SB_T2_WEST_SB_IN_B16_O)
	);
	corebit_and and_inst0(
		.in0(coreir_eq_16_inst0_out),
		.in1(config_read[0]),
		.out(and_inst0_out)
	);
	corebit_and and_inst1(
		.in0(coreir_eq_16_inst0_out),
		.in1(config_write[0]),
		.out(and_inst1_out)
	);
	coreir_const #(
		.value(8'h00),
		.width(8)
	) const_0_8(.out(const_0_8_out));
	coreir_const #(
		.value(9'h1ff),
		.width(9)
	) const_511_9(.out(const_511_9_out));
	coreir_eq #(.width(16)) coreir_eq_16_inst0(
		.in0(tile_id),
		.in1(self_config_config_addr_out[15:0]),
		.out(coreir_eq_16_inst0_out)
	);
	coreir_or #(.width(32)) read_config_data_or_inst0(
		.in0(read_data_mux_O),
		.in1(read_config_data_in),
		.out(read_config_data_or_inst0_out)
	);
	MuxWithDefaultWrapper_11_32_8_0 read_data_mux(
		.EN(and_inst0_out),
		.I_0(MemCore_inst0_read_config_data),
		.I_1(MemCore_inst0_read_config_data_1),
		.I_10(SB_ID0_3TRACKS_B16_MemCore_read_config_data),
		.I_2(CB_flush_read_config_data),
		.I_3(CB_input_width_16_num_0_read_config_data),
		.I_4(CB_input_width_16_num_1_read_config_data),
		.I_5(CB_input_width_16_num_2_read_config_data),
		.I_6(CB_input_width_16_num_3_read_config_data),
		.I_7(CB_input_width_1_num_0_read_config_data),
		.I_8(CB_input_width_1_num_1_read_config_data),
		.I_9(SB_ID0_3TRACKS_B1_MemCore_read_config_data),
		.O(read_data_mux_O),
		.S(read_data_mux_S_in)
	);
	mantle_wire__typeBitIn8 read_data_mux_S(
		.in(read_data_mux_S_in),
		.out(self_config_config_addr_out[23:16])
	);
	mantle_wire__typeBit32 self_config_config_addr(
		.in(config_config_addr),
		.out(self_config_config_addr_out)
	);
	assign SB_T0_EAST_SB_OUT_B1 = SB_ID0_3TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1;
	assign SB_T0_EAST_SB_OUT_B16 = SB_ID0_3TRACKS_B16_MemCore_SB_T0_EAST_SB_OUT_B16;
	assign SB_T0_NORTH_SB_OUT_B1 = SB_ID0_3TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1;
	assign SB_T0_NORTH_SB_OUT_B16 = SB_ID0_3TRACKS_B16_MemCore_SB_T0_NORTH_SB_OUT_B16;
	assign SB_T0_SOUTH_SB_OUT_B1 = SB_ID0_3TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1;
	assign SB_T0_SOUTH_SB_OUT_B16 = SB_ID0_3TRACKS_B16_MemCore_SB_T0_SOUTH_SB_OUT_B16;
	assign SB_T0_WEST_SB_OUT_B1 = SB_ID0_3TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1;
	assign SB_T0_WEST_SB_OUT_B16 = SB_ID0_3TRACKS_B16_MemCore_SB_T0_WEST_SB_OUT_B16;
	assign SB_T1_EAST_SB_OUT_B1 = SB_ID0_3TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1;
	assign SB_T1_EAST_SB_OUT_B16 = SB_ID0_3TRACKS_B16_MemCore_SB_T1_EAST_SB_OUT_B16;
	assign SB_T1_NORTH_SB_OUT_B1 = SB_ID0_3TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1;
	assign SB_T1_NORTH_SB_OUT_B16 = SB_ID0_3TRACKS_B16_MemCore_SB_T1_NORTH_SB_OUT_B16;
	assign SB_T1_SOUTH_SB_OUT_B1 = SB_ID0_3TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1;
	assign SB_T1_SOUTH_SB_OUT_B16 = SB_ID0_3TRACKS_B16_MemCore_SB_T1_SOUTH_SB_OUT_B16;
	assign SB_T1_WEST_SB_OUT_B1 = SB_ID0_3TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1;
	assign SB_T1_WEST_SB_OUT_B16 = SB_ID0_3TRACKS_B16_MemCore_SB_T1_WEST_SB_OUT_B16;
	assign SB_T2_EAST_SB_OUT_B1 = SB_ID0_3TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1;
	assign SB_T2_EAST_SB_OUT_B16 = SB_ID0_3TRACKS_B16_MemCore_SB_T2_EAST_SB_OUT_B16;
	assign SB_T2_NORTH_SB_OUT_B1 = SB_ID0_3TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1;
	assign SB_T2_NORTH_SB_OUT_B16 = SB_ID0_3TRACKS_B16_MemCore_SB_T2_NORTH_SB_OUT_B16;
	assign SB_T2_SOUTH_SB_OUT_B1 = SB_ID0_3TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1;
	assign SB_T2_SOUTH_SB_OUT_B16 = SB_ID0_3TRACKS_B16_MemCore_SB_T2_SOUTH_SB_OUT_B16;
	assign SB_T2_WEST_SB_OUT_B1 = SB_ID0_3TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1;
	assign SB_T2_WEST_SB_OUT_B16 = SB_ID0_3TRACKS_B16_MemCore_SB_T2_WEST_SB_OUT_B16;
	assign clk_out = clk_pass_through;
	assign clk_pass_through_out_bot = clk_pass_through;
	assign config_out_config_addr = config_config_addr;
	assign config_out_config_data = config_config_data;
	assign config_out_read = config_read;
	assign config_out_write = config_write;
	assign hi = const_511_9_out;
	assign lo = const_0_8_out;
	assign read_config_data = read_config_data_or_inst0_out;
	assign reset_out = reset;
	assign stall_out = stall;
endmodule
module CB_data1_sel (
	I,
	O
);
	input [3:0] I;
	output [3:0] O;
	assign O = I;
endmodule
module CB_data1 (
	I_0,
	I_1,
	I_10,
	I_11,
	I_2,
	I_3,
	I_4,
	I_5,
	I_6,
	I_7,
	I_8,
	I_9,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	read_config_data,
	reset
);
	input [15:0] I_0;
	input [15:0] I_1;
	input [15:0] I_10;
	input [15:0] I_11;
	input [15:0] I_2;
	input [15:0] I_3;
	input [15:0] I_4;
	input [15:0] I_5;
	input [15:0] I_6;
	input [15:0] I_7;
	input [15:0] I_8;
	input [15:0] I_9;
	output [15:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output [31:0] read_config_data;
	input reset;
	wire [3:0] CB_data1_sel_inst0_O;
	wire [15:0] MUX_CB_data1$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0_out;
	wire ZextWrapper_4_32_inst0$bit_const_0_None_out;
	wire [3:0] ZextWrapper_4_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_4_32_inst0$self_O_in;
	wire [3:0] config_reg_0_O;
	CB_data1_sel CB_data1_sel_inst0(
		.I(config_reg_0_O),
		.O(CB_data1_sel_inst0_O)
	);
	commonlib_muxn__N12__width16 MUX_CB_data1$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0(
		.in_data_0(I_0),
		.in_data_1(I_1),
		.in_data_10(I_10),
		.in_data_11(I_11),
		.in_data_2(I_2),
		.in_data_3(I_3),
		.in_data_4(I_4),
		.in_data_5(I_5),
		.in_data_6(I_6),
		.in_data_7(I_7),
		.in_data_8(I_8),
		.in_data_9(I_9),
		.in_sel(CB_data1_sel_inst0_O),
		.out(MUX_CB_data1$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_4_32_inst0$bit_const_0_None(.out(ZextWrapper_4_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit4 ZextWrapper_4_32_inst0$self_I(
		.in(config_reg_0_O),
		.out(ZextWrapper_4_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_4_32_inst0$self_O_out;
	assign ZextWrapper_4_32_inst0$self_O_out = {ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$self_I_out[3:0]};
	mantle_wire__typeBitIn32 ZextWrapper_4_32_inst0$self_O(
		.in(ZextWrapper_4_32_inst0$self_O_in),
		.out(ZextWrapper_4_32_inst0$self_O_out)
	);
	ConfigRegister_4_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = MUX_CB_data1$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0_out;
	assign read_config_data = ZextWrapper_4_32_inst0$self_O_in;
endmodule
module CB_data0_sel (
	I,
	O
);
	input [3:0] I;
	output [3:0] O;
	assign O = I;
endmodule
module CB_data0 (
	I_0,
	I_1,
	I_10,
	I_11,
	I_2,
	I_3,
	I_4,
	I_5,
	I_6,
	I_7,
	I_8,
	I_9,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	read_config_data,
	reset
);
	input [15:0] I_0;
	input [15:0] I_1;
	input [15:0] I_10;
	input [15:0] I_11;
	input [15:0] I_2;
	input [15:0] I_3;
	input [15:0] I_4;
	input [15:0] I_5;
	input [15:0] I_6;
	input [15:0] I_7;
	input [15:0] I_8;
	input [15:0] I_9;
	output [15:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output [31:0] read_config_data;
	input reset;
	wire [3:0] CB_data0_sel_inst0_O;
	wire [15:0] MUX_CB_data0$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0_out;
	wire ZextWrapper_4_32_inst0$bit_const_0_None_out;
	wire [3:0] ZextWrapper_4_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_4_32_inst0$self_O_in;
	wire [3:0] config_reg_0_O;
	CB_data0_sel CB_data0_sel_inst0(
		.I(config_reg_0_O),
		.O(CB_data0_sel_inst0_O)
	);
	commonlib_muxn__N12__width16 MUX_CB_data0$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0(
		.in_data_0(I_0),
		.in_data_1(I_1),
		.in_data_10(I_10),
		.in_data_11(I_11),
		.in_data_2(I_2),
		.in_data_3(I_3),
		.in_data_4(I_4),
		.in_data_5(I_5),
		.in_data_6(I_6),
		.in_data_7(I_7),
		.in_data_8(I_8),
		.in_data_9(I_9),
		.in_sel(CB_data0_sel_inst0_O),
		.out(MUX_CB_data0$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_4_32_inst0$bit_const_0_None(.out(ZextWrapper_4_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit4 ZextWrapper_4_32_inst0$self_I(
		.in(config_reg_0_O),
		.out(ZextWrapper_4_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_4_32_inst0$self_O_out;
	assign ZextWrapper_4_32_inst0$self_O_out = {ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$self_I_out[3:0]};
	mantle_wire__typeBitIn32 ZextWrapper_4_32_inst0$self_O(
		.in(ZextWrapper_4_32_inst0$self_O_in),
		.out(ZextWrapper_4_32_inst0$self_O_out)
	);
	ConfigRegister_4_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = MUX_CB_data0$Mux12xBits16_inst0$coreir_commonlib_mux12x16_inst0_out;
	assign read_config_data = ZextWrapper_4_32_inst0$self_O_in;
endmodule
module CB_bit2_sel (
	I,
	O
);
	input [3:0] I;
	output [3:0] O;
	assign O = I;
endmodule
module CB_bit2 (
	I_0,
	I_1,
	I_10,
	I_11,
	I_2,
	I_3,
	I_4,
	I_5,
	I_6,
	I_7,
	I_8,
	I_9,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	read_config_data,
	reset
);
	input [0:0] I_0;
	input [0:0] I_1;
	input [0:0] I_10;
	input [0:0] I_11;
	input [0:0] I_2;
	input [0:0] I_3;
	input [0:0] I_4;
	input [0:0] I_5;
	input [0:0] I_6;
	input [0:0] I_7;
	input [0:0] I_8;
	input [0:0] I_9;
	output [0:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output [31:0] read_config_data;
	input reset;
	wire [3:0] CB_bit2_sel_inst0_O;
	wire [0:0] MUX_CB_bit2$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0_out;
	wire ZextWrapper_4_32_inst0$bit_const_0_None_out;
	wire [3:0] ZextWrapper_4_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_4_32_inst0$self_O_in;
	wire [3:0] config_reg_0_O;
	CB_bit2_sel CB_bit2_sel_inst0(
		.I(config_reg_0_O),
		.O(CB_bit2_sel_inst0_O)
	);
	commonlib_muxn__N12__width1 MUX_CB_bit2$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0(
		.in_data_0(I_0),
		.in_data_1(I_1),
		.in_data_10(I_10),
		.in_data_11(I_11),
		.in_data_2(I_2),
		.in_data_3(I_3),
		.in_data_4(I_4),
		.in_data_5(I_5),
		.in_data_6(I_6),
		.in_data_7(I_7),
		.in_data_8(I_8),
		.in_data_9(I_9),
		.in_sel(CB_bit2_sel_inst0_O),
		.out(MUX_CB_bit2$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_4_32_inst0$bit_const_0_None(.out(ZextWrapper_4_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit4 ZextWrapper_4_32_inst0$self_I(
		.in(config_reg_0_O),
		.out(ZextWrapper_4_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_4_32_inst0$self_O_out;
	assign ZextWrapper_4_32_inst0$self_O_out = {ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$self_I_out[3:0]};
	mantle_wire__typeBitIn32 ZextWrapper_4_32_inst0$self_O(
		.in(ZextWrapper_4_32_inst0$self_O_in),
		.out(ZextWrapper_4_32_inst0$self_O_out)
	);
	ConfigRegister_4_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = MUX_CB_bit2$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0_out;
	assign read_config_data = ZextWrapper_4_32_inst0$self_O_in;
endmodule
module CB_bit1_sel (
	I,
	O
);
	input [3:0] I;
	output [3:0] O;
	assign O = I;
endmodule
module CB_bit1 (
	I_0,
	I_1,
	I_10,
	I_11,
	I_2,
	I_3,
	I_4,
	I_5,
	I_6,
	I_7,
	I_8,
	I_9,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	read_config_data,
	reset
);
	input [0:0] I_0;
	input [0:0] I_1;
	input [0:0] I_10;
	input [0:0] I_11;
	input [0:0] I_2;
	input [0:0] I_3;
	input [0:0] I_4;
	input [0:0] I_5;
	input [0:0] I_6;
	input [0:0] I_7;
	input [0:0] I_8;
	input [0:0] I_9;
	output [0:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output [31:0] read_config_data;
	input reset;
	wire [3:0] CB_bit1_sel_inst0_O;
	wire [0:0] MUX_CB_bit1$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0_out;
	wire ZextWrapper_4_32_inst0$bit_const_0_None_out;
	wire [3:0] ZextWrapper_4_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_4_32_inst0$self_O_in;
	wire [3:0] config_reg_0_O;
	CB_bit1_sel CB_bit1_sel_inst0(
		.I(config_reg_0_O),
		.O(CB_bit1_sel_inst0_O)
	);
	commonlib_muxn__N12__width1 MUX_CB_bit1$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0(
		.in_data_0(I_0),
		.in_data_1(I_1),
		.in_data_10(I_10),
		.in_data_11(I_11),
		.in_data_2(I_2),
		.in_data_3(I_3),
		.in_data_4(I_4),
		.in_data_5(I_5),
		.in_data_6(I_6),
		.in_data_7(I_7),
		.in_data_8(I_8),
		.in_data_9(I_9),
		.in_sel(CB_bit1_sel_inst0_O),
		.out(MUX_CB_bit1$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_4_32_inst0$bit_const_0_None(.out(ZextWrapper_4_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit4 ZextWrapper_4_32_inst0$self_I(
		.in(config_reg_0_O),
		.out(ZextWrapper_4_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_4_32_inst0$self_O_out;
	assign ZextWrapper_4_32_inst0$self_O_out = {ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$self_I_out[3:0]};
	mantle_wire__typeBitIn32 ZextWrapper_4_32_inst0$self_O(
		.in(ZextWrapper_4_32_inst0$self_O_in),
		.out(ZextWrapper_4_32_inst0$self_O_out)
	);
	ConfigRegister_4_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = MUX_CB_bit1$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0_out;
	assign read_config_data = ZextWrapper_4_32_inst0$self_O_in;
endmodule
module CB_bit0_sel (
	I,
	O
);
	input [3:0] I;
	output [3:0] O;
	assign O = I;
endmodule
module CB_bit0 (
	I_0,
	I_1,
	I_10,
	I_11,
	I_2,
	I_3,
	I_4,
	I_5,
	I_6,
	I_7,
	I_8,
	I_9,
	O,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	read_config_data,
	reset
);
	input [0:0] I_0;
	input [0:0] I_1;
	input [0:0] I_10;
	input [0:0] I_11;
	input [0:0] I_2;
	input [0:0] I_3;
	input [0:0] I_4;
	input [0:0] I_5;
	input [0:0] I_6;
	input [0:0] I_7;
	input [0:0] I_8;
	input [0:0] I_9;
	output [0:0] O;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	output [31:0] read_config_data;
	input reset;
	wire [3:0] CB_bit0_sel_inst0_O;
	wire [0:0] MUX_CB_bit0$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0_out;
	wire ZextWrapper_4_32_inst0$bit_const_0_None_out;
	wire [3:0] ZextWrapper_4_32_inst0$self_I_out;
	wire [31:0] ZextWrapper_4_32_inst0$self_O_in;
	wire [3:0] config_reg_0_O;
	CB_bit0_sel CB_bit0_sel_inst0(
		.I(config_reg_0_O),
		.O(CB_bit0_sel_inst0_O)
	);
	commonlib_muxn__N12__width1 MUX_CB_bit0$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0(
		.in_data_0(I_0),
		.in_data_1(I_1),
		.in_data_10(I_10),
		.in_data_11(I_11),
		.in_data_2(I_2),
		.in_data_3(I_3),
		.in_data_4(I_4),
		.in_data_5(I_5),
		.in_data_6(I_6),
		.in_data_7(I_7),
		.in_data_8(I_8),
		.in_data_9(I_9),
		.in_sel(CB_bit0_sel_inst0_O),
		.out(MUX_CB_bit0$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0_out)
	);
	corebit_const #(.value(1'b0)) ZextWrapper_4_32_inst0$bit_const_0_None(.out(ZextWrapper_4_32_inst0$bit_const_0_None_out));
	mantle_wire__typeBit4 ZextWrapper_4_32_inst0$self_I(
		.in(config_reg_0_O),
		.out(ZextWrapper_4_32_inst0$self_I_out)
	);
	wire [31:0] ZextWrapper_4_32_inst0$self_O_out;
	assign ZextWrapper_4_32_inst0$self_O_out = {ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$bit_const_0_None_out, ZextWrapper_4_32_inst0$self_I_out[3:0]};
	mantle_wire__typeBitIn32 ZextWrapper_4_32_inst0$self_O(
		.in(ZextWrapper_4_32_inst0$self_O_in),
		.out(ZextWrapper_4_32_inst0$self_O_out)
	);
	ConfigRegister_4_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	assign O = MUX_CB_bit0$Mux12xBits1_inst0$coreir_commonlib_mux12x1_inst0_out;
	assign read_config_data = ZextWrapper_4_32_inst0$self_O_in;
endmodule
module ALU (
	alu,
	signed_,
	a,
	b,
	d,
	O0,
	O1,
	O2,
	O3,
	O4,
	O5,
	CLK,
	ASYNCRESET
);
	input [7:0] alu;
	input [0:0] signed_;
	input [15:0] a;
	input [15:0] b;
	input d;
	output [15:0] O0;
	output O1;
	output O2;
	output O3;
	output O4;
	output O5;
	input CLK;
	input ASYNCRESET;
	wire [0:0] Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst13$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst14$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst15$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst16$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst17$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst18$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst19$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst20$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst21$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst22$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst23$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst24$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst25$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst26$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst27$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst28$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst29$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst30$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst31$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst32$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst33$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst34$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst35$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst36$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst37$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst38$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst39$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst40$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst41$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst42$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst43$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst44$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst45$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst46$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst47$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst48$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst49$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst50$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst51$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst52$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBit_inst9$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst10$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst11$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst12$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst13$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst14$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst15$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst16$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst17$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst18$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst18_I1_in;
	wire [15:0] Mux2xBits16_inst19$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst20$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst21$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst22$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst23$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst24$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst25$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst26$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst27$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst28$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst29$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst30$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst31$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst32$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst33$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst34$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst35$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst36$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst37$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst38$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst39$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst40$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst41$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst42$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst43$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst44$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst45$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst46$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst47$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst48$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst49$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst5$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst50$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst51$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst52$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst53$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst54$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst55$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst56$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst57$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst58$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst59$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst6$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst60$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst61$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst61_I1_in;
	wire [15:0] Mux2xBits16_inst62$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst63$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst64$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst64_I1_in;
	wire [15:0] Mux2xBits16_inst65$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst66$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst67$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst67_I1_in;
	wire [15:0] Mux2xBits16_inst68$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst69$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst70$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst70_I1_in;
	wire [15:0] Mux2xBits16_inst70_O_out;
	wire [15:0] Mux2xBits16_inst71$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst7_O_out;
	wire [15:0] Mux2xBits16_inst8$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xBits16_inst9$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [22:0] Mux2xBits23_inst0$coreir_commonlib_mux2x23_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst0$coreir_commonlib_mux2x8_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst0_I0_in;
	wire [7:0] Mux2xBits8_inst0_I1_in;
	wire [7:0] Mux2xBits8_inst1$coreir_commonlib_mux2x8_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst10$coreir_commonlib_mux2x8_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst10_I1_in;
	wire [7:0] Mux2xBits8_inst11$coreir_commonlib_mux2x8_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst11_I1_in;
	wire [7:0] Mux2xBits8_inst12$coreir_commonlib_mux2x8_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst12_I1_in;
	wire [7:0] Mux2xBits8_inst13$coreir_commonlib_mux2x8_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst13_I1_in;
	wire [7:0] Mux2xBits8_inst14$coreir_commonlib_mux2x8_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst14_I1_in;
	wire [7:0] Mux2xBits8_inst15$coreir_commonlib_mux2x8_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst15_I1_in;
	wire [7:0] Mux2xBits8_inst16$coreir_commonlib_mux2x8_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst16_I1_in;
	wire [7:0] Mux2xBits8_inst17$coreir_commonlib_mux2x8_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst17_I1_in;
	wire [7:0] Mux2xBits8_inst18$coreir_commonlib_mux2x8_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst18_I1_in;
	wire [7:0] Mux2xBits8_inst19$coreir_commonlib_mux2x8_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst19_I1_in;
	wire [7:0] Mux2xBits8_inst1_I1_in;
	wire [7:0] Mux2xBits8_inst2$coreir_commonlib_mux2x8_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst20$coreir_commonlib_mux2x8_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst20_I1_in;
	wire [7:0] Mux2xBits8_inst2_I1_in;
	wire [7:0] Mux2xBits8_inst3$coreir_commonlib_mux2x8_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst3_I1_in;
	wire [7:0] Mux2xBits8_inst4$coreir_commonlib_mux2x8_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst4_I1_in;
	wire [7:0] Mux2xBits8_inst5$coreir_commonlib_mux2x8_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst5_I1_in;
	wire [7:0] Mux2xBits8_inst6$coreir_commonlib_mux2x8_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst6_I1_in;
	wire [7:0] Mux2xBits8_inst7$coreir_commonlib_mux2x8_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst7_I1_in;
	wire [7:0] Mux2xBits8_inst8$coreir_commonlib_mux2x8_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst8_I1_in;
	wire [7:0] Mux2xBits8_inst9$coreir_commonlib_mux2x8_inst0$_join_out;
	wire [7:0] Mux2xBits8_inst9_I1_in;
	wire [15:0] Mux2xSInt16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst1$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst10$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst11$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst12$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst13$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst14$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst15$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst16$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst17$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst18$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst19$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst2$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst20$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst21$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst22$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst23$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst24$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst25$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst25_I1_in;
	wire [15:0] Mux2xSInt16_inst26$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst27$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst28$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst28_I0_in;
	wire [15:0] Mux2xSInt16_inst29$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst3$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst30$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst4$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst5$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst6$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst7$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [15:0] Mux2xSInt16_inst9$coreir_commonlib_mux2x16_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst0$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst0_O_out;
	wire [8:0] Mux2xSInt9_inst1$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst10$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst11$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst11_I1_in;
	wire [8:0] Mux2xSInt9_inst12$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst13$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst13_I1_in;
	wire [8:0] Mux2xSInt9_inst14$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst15$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst15_I1_in;
	wire [8:0] Mux2xSInt9_inst16$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst17$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst17_I1_in;
	wire [8:0] Mux2xSInt9_inst18$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst19$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst19_I1_in;
	wire [8:0] Mux2xSInt9_inst1_I0_in;
	wire [8:0] Mux2xSInt9_inst1_I1_in;
	wire [8:0] Mux2xSInt9_inst2$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst20$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst21$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst21_I1_in;
	wire [8:0] Mux2xSInt9_inst22$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst23$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst23_I1_in;
	wire [8:0] Mux2xSInt9_inst24$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst25$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst25_I1_in;
	wire [8:0] Mux2xSInt9_inst26$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst27$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst27_I1_in;
	wire [8:0] Mux2xSInt9_inst28$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst29$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst29_I1_in;
	wire [8:0] Mux2xSInt9_inst3$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst30$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst31$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst31_I1_in;
	wire [8:0] Mux2xSInt9_inst32$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst33$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst33_I1_in;
	wire [8:0] Mux2xSInt9_inst34$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst35$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst35_I1_in;
	wire [8:0] Mux2xSInt9_inst36$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst37$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst37_I1_in;
	wire [8:0] Mux2xSInt9_inst38$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst39$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst39_I1_in;
	wire [8:0] Mux2xSInt9_inst3_I1_in;
	wire [8:0] Mux2xSInt9_inst4$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst40$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst41$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst41_I1_in;
	wire [8:0] Mux2xSInt9_inst42$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst5$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst5_I1_in;
	wire [8:0] Mux2xSInt9_inst6$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst7$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst7_I1_in;
	wire [8:0] Mux2xSInt9_inst8$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst9$coreir_commonlib_mux2x9_inst0$_join_out;
	wire [8:0] Mux2xSInt9_inst9_I1_in;
	wire [31:0] Mux2xUInt32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
	wire [31:0] Mux2xUInt32_inst0_I0_in;
	wire [31:0] Mux2xUInt32_inst0_I1_in;
	wire [31:0] Mux2xUInt32_inst1$coreir_commonlib_mux2x32_inst0$_join_out;
	wire [31:0] Mux2xUInt32_inst1_I0_in;
	wire [31:0] Mux2xUInt32_inst1_I1_in;
	wire bit_const_0_None_out;
	wire bit_const_1_None_out;
	wire [15:0] const_0_16_out;
	wire [22:0] const_0_23_out;
	wire [6:0] const_0_7_out;
	wire [7:0] const_0_8_out;
	wire [8:0] const_0_9_out;
	wire [15:0] const_10_16_out;
	wire [15:0] const_11_16_out;
	wire [7:0] const_11_8_out;
	wire [15:0] const_127_16_out;
	wire [7:0] const_127_8_out;
	wire [8:0] const_127_9_out;
	wire [15:0] const_128_16_out;
	wire [15:0] const_12_16_out;
	wire [7:0] const_12_8_out;
	wire [15:0] const_13_16_out;
	wire [7:0] const_13_8_out;
	wire [7:0] const_142_8_out;
	wire [7:0] const_146_8_out;
	wire [7:0] const_147_8_out;
	wire [7:0] const_148_8_out;
	wire [7:0] const_149_8_out;
	wire [15:0] const_14_16_out;
	wire [7:0] const_150_8_out;
	wire [7:0] const_151_8_out;
	wire [7:0] const_152_8_out;
	wire [15:0] const_15_16_out;
	wire [7:0] const_15_8_out;
	wire [7:0] const_17_8_out;
	wire [7:0] const_18_8_out;
	wire [7:0] const_19_8_out;
	wire [0:0] const_1_1_out;
	wire [15:0] const_1_16_out;
	wire [7:0] const_1_8_out;
	wire [7:0] const_20_8_out;
	wire [7:0] const_22_8_out;
	wire [7:0] const_23_8_out;
	wire [7:0] const_24_8_out;
	wire [7:0] const_255_8_out;
	wire [8:0] const_255_9_out;
	wire [7:0] const_25_8_out;
	wire [15:0] const_2_16_out;
	wire [7:0] const_2_8_out;
	wire [15:0] const_32512_16_out;
	wire [15:0] const_32640_16_out;
	wire [15:0] const_32768_16_out;
	wire [15:0] const_3_16_out;
	wire [7:0] const_3_8_out;
	wire [15:0] const_4_16_out;
	wire [7:0] const_4_8_out;
	wire [15:0] const_5_16_out;
	wire [7:0] const_5_8_out;
	wire [15:0] const_65409_16_out;
	wire [15:0] const_6_16_out;
	wire [7:0] const_6_8_out;
	wire [15:0] const_7_16_out;
	wire [22:0] const_7_23_out;
	wire [15:0] const_8_16_out;
	wire [7:0] const_8_8_out;
	wire [15:0] const_9_16_out;
	wire [15:0] magma_BFloat_16_add_inst0_out;
	wire [15:0] magma_BFloat_16_mul_inst0_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bit_and_inst1_out;
	wire magma_Bit_and_inst2_out;
	wire magma_Bit_and_inst3_out;
	wire magma_Bit_and_inst4_out;
	wire magma_Bit_and_inst5_out;
	wire magma_Bit_and_inst6_out;
	wire magma_Bit_and_inst7_out;
	wire magma_Bit_and_inst8_out;
	wire magma_Bit_not_inst0_out;
	wire magma_Bit_not_inst1_out;
	wire magma_Bit_not_inst10_out;
	wire magma_Bit_not_inst11_out;
	wire magma_Bit_not_inst12_out;
	wire magma_Bit_not_inst13_out;
	wire magma_Bit_not_inst14_out;
	wire magma_Bit_not_inst15_out;
	wire magma_Bit_not_inst16_out;
	wire magma_Bit_not_inst17_out;
	wire magma_Bit_not_inst18_out;
	wire magma_Bit_not_inst19_out;
	wire magma_Bit_not_inst2_out;
	wire magma_Bit_not_inst20_out;
	wire magma_Bit_not_inst21_out;
	wire magma_Bit_not_inst22_out;
	wire magma_Bit_not_inst23_out;
	wire magma_Bit_not_inst24_out;
	wire magma_Bit_not_inst25_out;
	wire magma_Bit_not_inst26_out;
	wire magma_Bit_not_inst27_out;
	wire magma_Bit_not_inst28_out;
	wire magma_Bit_not_inst3_out;
	wire magma_Bit_not_inst4_out;
	wire magma_Bit_not_inst5_out;
	wire magma_Bit_not_inst6_out;
	wire magma_Bit_not_inst7_out;
	wire magma_Bit_not_inst8_out;
	wire magma_Bit_not_inst9_out;
	wire magma_Bit_or_inst0_out;
	wire magma_Bit_or_inst1_out;
	wire magma_Bit_or_inst10_out;
	wire magma_Bit_or_inst11_out;
	wire magma_Bit_or_inst12_out;
	wire magma_Bit_or_inst13_out;
	wire magma_Bit_or_inst2_out;
	wire magma_Bit_or_inst3_out;
	wire magma_Bit_or_inst4_out;
	wire magma_Bit_or_inst5_out;
	wire magma_Bit_or_inst6_out;
	wire magma_Bit_or_inst7_out;
	wire magma_Bit_or_inst8_out;
	wire magma_Bit_or_inst9_out;
	wire magma_Bit_xor_inst0_out;
	wire magma_Bit_xor_inst1_out;
	wire magma_Bit_xor_inst10_out;
	wire magma_Bit_xor_inst11_out;
	wire magma_Bit_xor_inst12_out;
	wire magma_Bit_xor_inst13_out;
	wire magma_Bit_xor_inst14_out;
	wire magma_Bit_xor_inst15_out;
	wire magma_Bit_xor_inst16_out;
	wire magma_Bit_xor_inst17_out;
	wire magma_Bit_xor_inst18_out;
	wire magma_Bit_xor_inst19_out;
	wire magma_Bit_xor_inst2_out;
	wire magma_Bit_xor_inst20_out;
	wire magma_Bit_xor_inst21_out;
	wire magma_Bit_xor_inst22_out;
	wire magma_Bit_xor_inst23_out;
	wire magma_Bit_xor_inst24_out;
	wire magma_Bit_xor_inst25_out;
	wire magma_Bit_xor_inst3_out;
	wire magma_Bit_xor_inst4_out;
	wire magma_Bit_xor_inst5_out;
	wire magma_Bit_xor_inst6_out;
	wire magma_Bit_xor_inst7_out;
	wire magma_Bit_xor_inst8_out;
	wire magma_Bit_xor_inst9_out;
	wire [15:0] magma_Bits_16_and_inst0_out;
	wire [15:0] magma_Bits_16_and_inst1_out;
	wire [15:0] magma_Bits_16_and_inst10_out;
	wire [15:0] magma_Bits_16_and_inst11_out;
	wire [15:0] magma_Bits_16_and_inst12_out;
	wire [15:0] magma_Bits_16_and_inst13_out;
	wire [15:0] magma_Bits_16_and_inst14_out;
	wire [15:0] magma_Bits_16_and_inst15_out;
	wire [15:0] magma_Bits_16_and_inst16_out;
	wire [15:0] magma_Bits_16_and_inst17_out;
	wire [15:0] magma_Bits_16_and_inst2_out;
	wire [15:0] magma_Bits_16_and_inst3_out;
	wire [15:0] magma_Bits_16_and_inst4_out;
	wire [15:0] magma_Bits_16_and_inst5_out;
	wire [15:0] magma_Bits_16_and_inst6_out;
	wire [15:0] magma_Bits_16_and_inst7_out;
	wire [15:0] magma_Bits_16_and_inst8_out;
	wire [15:0] magma_Bits_16_and_inst9_out;
	wire magma_Bits_16_eq_inst0_out;
	wire magma_Bits_16_eq_inst1_out;
	wire [15:0] magma_Bits_16_lshr_inst0_out;
	wire [15:0] magma_Bits_16_lshr_inst1_out;
	wire [15:0] magma_Bits_16_not_inst0_out;
	wire [15:0] magma_Bits_16_or_inst0_out;
	wire [15:0] magma_Bits_16_or_inst1_out;
	wire [15:0] magma_Bits_16_or_inst2_out;
	wire [15:0] magma_Bits_16_or_inst3_out;
	wire [15:0] magma_Bits_16_or_inst4_out;
	wire [15:0] magma_Bits_16_or_inst5_out;
	wire [15:0] magma_Bits_16_or_inst6_out;
	wire [15:0] magma_Bits_16_or_inst7_out;
	wire [15:0] magma_Bits_16_or_inst8_out;
	wire [15:0] magma_Bits_16_or_inst9_out;
	wire [15:0] magma_Bits_16_shl_inst0_out;
	wire [15:0] magma_Bits_16_shl_inst1_out;
	wire [15:0] magma_Bits_16_shl_inst2_out;
	wire [15:0] magma_Bits_16_shl_inst3_out;
	wire [15:0] magma_Bits_16_shl_inst4_out;
	wire [15:0] magma_Bits_16_shl_inst5_out;
	wire [15:0] magma_Bits_16_xor_inst0_out;
	wire [15:0] magma_Bits_16_xor_inst1_out;
	wire magma_Bits_1_eq_inst0_out;
	wire magma_Bits_1_eq_inst1_out;
	wire [22:0] magma_Bits_23_lshr_inst0_out;
	wire [22:0] magma_Bits_23_shl_inst0_out;
	wire magma_Bits_7_eq_inst0_out;
	wire magma_Bits_7_eq_inst1_out;
	wire magma_Bits_7_eq_inst2_out;
	wire magma_Bits_8_eq_inst0_out;
	wire magma_Bits_8_eq_inst1_out;
	wire magma_Bits_8_eq_inst10_out;
	wire magma_Bits_8_eq_inst11_out;
	wire magma_Bits_8_eq_inst12_out;
	wire magma_Bits_8_eq_inst13_out;
	wire magma_Bits_8_eq_inst14_out;
	wire magma_Bits_8_eq_inst15_out;
	wire magma_Bits_8_eq_inst16_out;
	wire magma_Bits_8_eq_inst17_out;
	wire magma_Bits_8_eq_inst18_out;
	wire magma_Bits_8_eq_inst19_out;
	wire magma_Bits_8_eq_inst2_out;
	wire magma_Bits_8_eq_inst20_out;
	wire magma_Bits_8_eq_inst21_out;
	wire magma_Bits_8_eq_inst22_out;
	wire magma_Bits_8_eq_inst23_out;
	wire magma_Bits_8_eq_inst24_out;
	wire magma_Bits_8_eq_inst25_out;
	wire magma_Bits_8_eq_inst26_out;
	wire magma_Bits_8_eq_inst27_out;
	wire magma_Bits_8_eq_inst28_out;
	wire magma_Bits_8_eq_inst29_out;
	wire magma_Bits_8_eq_inst3_out;
	wire magma_Bits_8_eq_inst30_out;
	wire magma_Bits_8_eq_inst31_out;
	wire magma_Bits_8_eq_inst32_out;
	wire magma_Bits_8_eq_inst33_out;
	wire magma_Bits_8_eq_inst34_out;
	wire magma_Bits_8_eq_inst35_out;
	wire magma_Bits_8_eq_inst36_out;
	wire magma_Bits_8_eq_inst37_out;
	wire magma_Bits_8_eq_inst38_out;
	wire magma_Bits_8_eq_inst39_out;
	wire magma_Bits_8_eq_inst4_out;
	wire magma_Bits_8_eq_inst40_out;
	wire magma_Bits_8_eq_inst41_out;
	wire magma_Bits_8_eq_inst42_out;
	wire magma_Bits_8_eq_inst5_out;
	wire magma_Bits_8_eq_inst6_out;
	wire magma_Bits_8_eq_inst7_out;
	wire magma_Bits_8_eq_inst8_out;
	wire magma_Bits_8_eq_inst9_out;
	wire [15:0] magma_SInt_16_add_inst0_out;
	wire [15:0] magma_SInt_16_and_inst0_out;
	wire [15:0] magma_SInt_16_ashr_inst0_out;
	wire magma_SInt_16_eq_inst0_out;
	wire [15:0] magma_SInt_16_neg_inst0_out;
	wire [15:0] magma_SInt_16_neg_inst1_out;
	wire [15:0] magma_SInt_16_neg_inst2_out;
	wire [15:0] magma_SInt_16_neg_inst3_out;
	wire magma_SInt_16_sge_inst0_out;
	wire magma_SInt_16_sge_inst1_out;
	wire magma_SInt_16_sge_inst2_out;
	wire [15:0] magma_SInt_16_shl_inst0_out;
	wire magma_SInt_16_sle_inst0_out;
	wire [15:0] magma_SInt_16_sub_inst0_out;
	wire [15:0] magma_SInt_16_sub_inst1_out;
	wire [8:0] magma_SInt_9_neg_inst0_out;
	wire [8:0] magma_SInt_9_neg_inst1_out;
	wire magma_SInt_9_slt_inst0_out;
	wire magma_SInt_9_slt_inst1_out;
	wire magma_SInt_9_slt_inst2_out;
	wire [8:0] magma_SInt_9_sub_inst0_out;
	wire [8:0] magma_SInt_9_sub_inst1_out;
	wire [8:0] magma_SInt_9_sub_inst2_out;
	wire [15:0] magma_UInt_16_lshr_inst0_out;
	wire magma_UInt_16_uge_inst0_out;
	wire magma_UInt_16_ule_inst0_out;
	wire [16:0] magma_UInt_17_add_inst0_out;
	wire [16:0] magma_UInt_17_add_inst1_out;
	wire [31:0] magma_UInt_32_and_inst0_out;
	wire [31:0] magma_UInt_32_and_inst1_out;
	wire [31:0] magma_UInt_32_mul_inst0_out;
	wire [7:0] magma_UInt_8_add_inst0_out;
	wire [7:0] magma_UInt_8_add_inst1_out;
	wire [7:0] magma_UInt_8_sub_inst0_out;
	wire magma_UInt_8_ugt_inst0_out;
	wire [8:0] magma_UInt_9_add_inst0_out;
	wire magma_UInt_9_ugt_inst0_out;
	coreir_mux #(.width(1)) Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(bit_const_1_None_out),
		.in1(magma_SInt_16_sge_inst1_out),
		.sel(magma_Bits_1_eq_inst0_out),
		.out(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join(
		.in0(magma_UInt_16_uge_inst0_out),
		.in1(magma_SInt_16_sge_inst0_out),
		.sel(magma_Bits_1_eq_inst0_out),
		.out(Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst10$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst33_out),
		.out(Mux2xBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst11$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst9$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst33_out),
		.out(Mux2xBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst12$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst32_out),
		.out(Mux2xBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst13$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(magma_UInt_9_ugt_inst0_out),
		.sel(magma_Bits_8_eq_inst32_out),
		.out(Mux2xBit_inst13$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst14$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst31_out),
		.out(Mux2xBit_inst14$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst15$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst13$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst31_out),
		.out(Mux2xBit_inst15$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst16$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst14$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst30_out),
		.out(Mux2xBit_inst16$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst17$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst15$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst30_out),
		.out(Mux2xBit_inst17$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst18$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst16$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bit_or_inst7_out),
		.out(Mux2xBit_inst18$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst19$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst17$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bit_or_inst7_out),
		.out(Mux2xBit_inst19$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join(
		.in0(magma_UInt_16_ule_inst0_out),
		.in1(magma_SInt_16_sle_inst0_out),
		.sel(magma_Bits_1_eq_inst0_out),
		.out(Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst20$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst18$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst24_out),
		.out(Mux2xBit_inst20$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst21$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst19$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst24_out),
		.out(Mux2xBit_inst21$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst22$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst20$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst23_out),
		.out(Mux2xBit_inst22$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst23$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst21$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst23_out),
		.out(Mux2xBit_inst23$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst24$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst22$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst22_out),
		.out(Mux2xBit_inst24$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst25$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst23$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst22_out),
		.out(Mux2xBit_inst25$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst26$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst24$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst21_out),
		.out(Mux2xBit_inst26$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst27$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst25$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst21_out),
		.out(Mux2xBit_inst27$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst28$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst26$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst20_out),
		.out(Mux2xBit_inst28$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst29$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst27$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst20_out),
		.out(Mux2xBit_inst29$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join(
		.in0(bit_const_0_None_out),
		.in1(d),
		.sel(magma_Bit_or_inst1_out),
		.out(Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst30$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst28$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst19_out),
		.out(Mux2xBit_inst30$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst31$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst29$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst19_out),
		.out(Mux2xBit_inst31$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst32$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst30$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst18_out),
		.out(Mux2xBit_inst32$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst33$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst31$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(a[15]),
		.sel(magma_Bits_8_eq_inst18_out),
		.out(Mux2xBit_inst33$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst34$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst32$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst17_out),
		.out(Mux2xBit_inst34$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst35$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst33$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.sel(magma_Bits_8_eq_inst17_out),
		.out(Mux2xBit_inst35$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst36$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst34$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst16_out),
		.out(Mux2xBit_inst36$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst37$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst35$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.sel(magma_Bits_8_eq_inst16_out),
		.out(Mux2xBit_inst37$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst38$coreir_commonlib_mux2x1_inst0$_join(
		.in0(bit_const_0_None_out),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst15_out),
		.out(Mux2xBit_inst38$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst39$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst36$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst15_out),
		.out(Mux2xBit_inst39$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_1_None_out),
		.sel(magma_Bits_8_eq_inst6_out),
		.out(Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst40$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst37$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst15_out),
		.out(Mux2xBit_inst40$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst41$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst38$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst14_out),
		.out(Mux2xBit_inst41$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst42$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst39$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst14_out),
		.out(Mux2xBit_inst42$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst43$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst40$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst14_out),
		.out(Mux2xBit_inst43$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst44$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst41$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst13_out),
		.out(Mux2xBit_inst44$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst45$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst42$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst13_out),
		.out(Mux2xBit_inst45$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst46$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst43$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst13_out),
		.out(Mux2xBit_inst46$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst47$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst44$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(magma_UInt_17_add_inst1_out[16]),
		.sel(magma_Bit_or_inst4_out),
		.out(Mux2xBit_inst47$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst48$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst45$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(magma_Bit_or_inst5_out),
		.sel(magma_Bit_or_inst4_out),
		.out(Mux2xBit_inst48$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst49$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst46$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(magma_UInt_17_add_inst1_out[16]),
		.sel(magma_Bit_or_inst4_out),
		.out(Mux2xBit_inst49$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst5$coreir_commonlib_mux2x1_inst0$_join(
		.in0(bit_const_0_None_out),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst36_out),
		.out(Mux2xBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst50$coreir_commonlib_mux2x1_inst0$_join(
		.in0(magma_SInt_16_eq_inst0_out),
		.in1(magma_Bit_and_inst6_out),
		.sel(magma_Bit_or_inst11_out),
		.out(Mux2xBit_inst50$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst51$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst50$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_1_None_out),
		.sel(magma_Bit_and_inst8_out),
		.out(Mux2xBit_inst51$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst52$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst50$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(Mux2xBit_inst51$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.sel(magma_Bits_8_eq_inst42_out),
		.out(Mux2xBit_inst52$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst6$coreir_commonlib_mux2x1_inst0$_join(
		.in0(bit_const_0_None_out),
		.in1(magma_UInt_8_ugt_inst0_out),
		.sel(magma_Bits_8_eq_inst35_out),
		.out(Mux2xBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst7$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst35_out),
		.out(Mux2xBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst8$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst34_out),
		.out(Mux2xBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBit_inst9$coreir_commonlib_mux2x1_inst0$_join(
		.in0(Mux2xBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.in1(bit_const_0_None_out),
		.sel(magma_Bits_8_eq_inst34_out),
		.out(Mux2xBit_inst9$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(magma_UInt_16_lshr_inst0_out),
		.in1(magma_SInt_16_ashr_inst0_out),
		.sel(magma_Bits_1_eq_inst0_out),
		.out(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join(
		.in0(const_0_16_out),
		.in1(const_32768_16_out),
		.sel(magma_SInt_9_slt_inst0_out),
		.out(Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst10$coreir_commonlib_mux2x16_inst0$_join(
		.in0(magma_SInt_16_neg_inst1_out),
		.in1(a),
		.sel(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.out(Mux2xBits16_inst10$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst11$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(a),
		.sel(d),
		.out(Mux2xBits16_inst11$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst12$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(magma_Bits_16_xor_inst1_out),
		.sel(magma_Bit_or_inst8_out),
		.out(Mux2xBits16_inst12$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst13$coreir_commonlib_mux2x16_inst0$_join(
		.in0(magma_Bits_16_shl_inst5_out),
		.in1(magma_Bits_16_lshr_inst1_out),
		.sel(magma_SInt_9_slt_inst2_out),
		.out(Mux2xBits16_inst13$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst14$coreir_commonlib_mux2x16_inst0$_join(
		.in0(magma_Bits_16_or_inst1_out),
		.in1(Mux2xSInt16_inst29$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst36_out),
		.out(Mux2xBits16_inst14$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst15$coreir_commonlib_mux2x16_inst0$_join(
		.in0(magma_Bits_16_or_inst9_out),
		.in1(magma_Bits_16_or_inst8_out),
		.sel(magma_Bits_8_eq_inst35_out),
		.out(Mux2xBits16_inst15$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst16$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst14$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xSInt16_inst28$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst35_out),
		.out(Mux2xBits16_inst16$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst17$coreir_commonlib_mux2x16_inst0$_join(
		.in0(magma_Bits_16_and_inst11_out),
		.in1(magma_Bits_16_and_inst9_out),
		.sel(magma_Bits_8_eq_inst35_out),
		.out(Mux2xBits16_inst17$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst18$coreir_commonlib_mux2x16_inst0$_join(
		.in0(magma_Bits_16_and_inst13_out),
		.in1(Mux2xBits16_inst18_I1_in),
		.sel(magma_Bits_8_eq_inst35_out),
		.out(Mux2xBits16_inst18$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	mantle_wire__typeBitIn16 Mux2xBits16_inst18_I1(
		.in(Mux2xBits16_inst18_I1_in),
		.out(magma_Bits_23_lshr_inst0_out[15:0])
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst19$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst16$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(magma_Bits_16_or_inst1_out),
		.sel(magma_Bits_8_eq_inst34_out),
		.out(Mux2xBits16_inst19$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join(
		.in0(const_0_16_out),
		.in1(magma_Bits_16_and_inst0_out),
		.sel(magma_Bits_1_eq_inst1_out),
		.out(Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst20$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst15$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(magma_Bits_16_and_inst8_out),
		.sel(magma_Bits_8_eq_inst33_out),
		.out(Mux2xBits16_inst20$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst21$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst19$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(magma_Bits_16_or_inst7_out),
		.sel(magma_Bits_8_eq_inst33_out),
		.out(Mux2xBits16_inst21$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst22$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst17$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(magma_Bits_16_and_inst6_out),
		.sel(magma_Bits_8_eq_inst33_out),
		.out(Mux2xBits16_inst22$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst23$coreir_commonlib_mux2x16_inst0$_join(
		.in0(magma_Bits_16_shl_inst4_out),
		.in1(magma_Bits_16_shl_inst3_out),
		.sel(magma_Bits_8_eq_inst32_out),
		.out(Mux2xBits16_inst23$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst24$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst21$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(magma_Bits_16_or_inst4_out),
		.sel(magma_Bits_8_eq_inst32_out),
		.out(Mux2xBits16_inst24$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst25$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(magma_Bits_16_and_inst4_out),
		.sel(magma_Bits_8_eq_inst32_out),
		.out(Mux2xBits16_inst25$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst26$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst24$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(magma_Bits_16_and_inst3_out),
		.sel(magma_Bits_8_eq_inst31_out),
		.out(Mux2xBits16_inst26$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst27$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst25$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst31_out),
		.out(Mux2xBits16_inst27$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst28$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst26$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(magma_BFloat_16_mul_inst0_out),
		.sel(magma_Bits_8_eq_inst30_out),
		.out(Mux2xBits16_inst28$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst29$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst27$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst30_out),
		.out(Mux2xBits16_inst29$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join(
		.in0(a),
		.in1(magma_SInt_16_neg_inst0_out),
		.sel(magma_Bit_not_inst8_out),
		.out(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst30$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst12$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bit_or_inst7_out),
		.out(Mux2xBits16_inst30$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst31$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst28$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(magma_BFloat_16_add_inst0_out),
		.sel(magma_Bit_or_inst7_out),
		.out(Mux2xBits16_inst31$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst32$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst29$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bit_or_inst7_out),
		.out(Mux2xBits16_inst32$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst33$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst30$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst24_out),
		.out(Mux2xBits16_inst33$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst34$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst31$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(magma_Bits_16_shl_inst1_out),
		.sel(magma_Bits_8_eq_inst24_out),
		.out(Mux2xBits16_inst34$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst35$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst32$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst24_out),
		.out(Mux2xBits16_inst35$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst36$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst33$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst23_out),
		.out(Mux2xBits16_inst36$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst37$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst34$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst23_out),
		.out(Mux2xBits16_inst37$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst38$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst35$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst23_out),
		.out(Mux2xBits16_inst38$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst39$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst36$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst22_out),
		.out(Mux2xBits16_inst39$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst2_out),
		.out(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst40$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst37$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(magma_Bits_16_xor_inst0_out),
		.sel(magma_Bits_8_eq_inst22_out),
		.out(Mux2xBits16_inst40$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst41$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst38$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst22_out),
		.out(Mux2xBits16_inst41$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst42$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst39$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst21_out),
		.out(Mux2xBits16_inst42$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst43$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst40$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(magma_Bits_16_or_inst2_out),
		.sel(magma_Bits_8_eq_inst21_out),
		.out(Mux2xBits16_inst43$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst44$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst41$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst21_out),
		.out(Mux2xBits16_inst44$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst45$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst42$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst20_out),
		.out(Mux2xBits16_inst45$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst46$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst43$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(magma_Bits_16_and_inst2_out),
		.sel(magma_Bits_8_eq_inst20_out),
		.out(Mux2xBits16_inst46$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst47$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst44$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst20_out),
		.out(Mux2xBits16_inst47$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst48$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst45$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst19_out),
		.out(Mux2xBits16_inst48$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst49$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst46$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst11$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst19_out),
		.out(Mux2xBits16_inst49$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst5$coreir_commonlib_mux2x16_inst0$_join(
		.in0(const_0_16_out),
		.in1(magma_SInt_16_and_inst0_out),
		.sel(magma_SInt_16_sge_inst2_out),
		.out(Mux2xBits16_inst5$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst50$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst47$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst19_out),
		.out(Mux2xBits16_inst50$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst51$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst48$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst18_out),
		.out(Mux2xBits16_inst51$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst52$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst49$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst10$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst18_out),
		.out(Mux2xBits16_inst52$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst53$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst50$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst18_out),
		.out(Mux2xBits16_inst53$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst54$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst51$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst17_out),
		.out(Mux2xBits16_inst54$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst55$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst52$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst9$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst17_out),
		.out(Mux2xBits16_inst55$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst56$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst53$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst17_out),
		.out(Mux2xBits16_inst56$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst57$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst54$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst16_out),
		.out(Mux2xBits16_inst57$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst58$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst55$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst8$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst16_out),
		.out(Mux2xBits16_inst58$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst59$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst56$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst16_out),
		.out(Mux2xBits16_inst59$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst6$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst5$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(magma_Bits_16_lshr_inst0_out),
		.sel(magma_Bits_8_eq_inst3_out),
		.out(Mux2xBits16_inst6$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst60$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst57$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst15_out),
		.out(Mux2xBits16_inst60$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst61$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst58$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst61_I1_in),
		.sel(magma_Bits_8_eq_inst15_out),
		.out(Mux2xBits16_inst61$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	mantle_wire__typeBitIn16 Mux2xBits16_inst61_I1(
		.in(Mux2xBits16_inst61_I1_in),
		.out(magma_UInt_32_mul_inst0_out[31:16])
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst62$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst59$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst15_out),
		.out(Mux2xBits16_inst62$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst63$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst60$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst14_out),
		.out(Mux2xBits16_inst63$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst64$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst61$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst64_I1_in),
		.sel(magma_Bits_8_eq_inst14_out),
		.out(Mux2xBits16_inst64$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	mantle_wire__typeBitIn16 Mux2xBits16_inst64_I1(
		.in(Mux2xBits16_inst64_I1_in),
		.out(magma_UInt_32_mul_inst0_out[23:8])
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst65$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst62$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst14_out),
		.out(Mux2xBits16_inst65$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst66$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst63$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst13_out),
		.out(Mux2xBits16_inst66$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst67$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst64$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst67_I1_in),
		.sel(magma_Bits_8_eq_inst13_out),
		.out(Mux2xBits16_inst67$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	mantle_wire__typeBitIn16 Mux2xBits16_inst67_I1(
		.in(Mux2xBits16_inst67_I1_in),
		.out(magma_UInt_32_mul_inst0_out[15:0])
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst68$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst65$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst13_out),
		.out(Mux2xBits16_inst68$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst69$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst66$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bit_or_inst4_out),
		.out(Mux2xBits16_inst69$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join(
		.in0(b),
		.in1(magma_Bits_16_not_inst0_out),
		.sel(magma_Bit_or_inst0_out),
		.out(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst70$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst67$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst70_I1_in),
		.sel(magma_Bit_or_inst4_out),
		.out(Mux2xBits16_inst70$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	mantle_wire__typeBitIn16 Mux2xBits16_inst70_I1(
		.in(Mux2xBits16_inst70_I1_in),
		.out(magma_UInt_17_add_inst1_out[15:0])
	);
	mantle_wire__typeBit16 Mux2xBits16_inst70_O(
		.in(Mux2xBits16_inst70$coreir_commonlib_mux2x16_inst0$_join_out),
		.out(Mux2xBits16_inst70_O_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst71$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst68$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bit_or_inst4_out),
		.out(Mux2xBits16_inst71$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	mantle_wire__typeBit16 Mux2xBits16_inst7_O(
		.in(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.out(Mux2xBits16_inst7_O_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst8$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(a),
		.sel(Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.out(Mux2xBits16_inst8$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xBits16_inst9$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(a),
		.sel(Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out[0]),
		.out(Mux2xBits16_inst9$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(23)) Mux2xBits23_inst0$coreir_commonlib_mux2x23_inst0$_join(
		.in0(magma_Bits_23_shl_inst0_out),
		.in1(const_0_23_out),
		.sel(magma_SInt_9_slt_inst1_out),
		.out(Mux2xBits23_inst0$coreir_commonlib_mux2x23_inst0$_join_out)
	);
	coreir_mux #(.width(8)) Mux2xBits8_inst0$coreir_commonlib_mux2x8_inst0$_join(
		.in0(Mux2xBits8_inst0_I0_in),
		.in1(Mux2xBits8_inst0_I1_in),
		.sel(magma_Bits_8_eq_inst36_out),
		.out(Mux2xBits8_inst0$coreir_commonlib_mux2x8_inst0$_join_out)
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst0_I0(
		.in(Mux2xBits8_inst0_I0_in),
		.out(a[14:7])
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst0_I1(
		.in(Mux2xBits8_inst0_I1_in),
		.out(a[14:7])
	);
	coreir_mux #(.width(8)) Mux2xBits8_inst1$coreir_commonlib_mux2x8_inst0$_join(
		.in0(Mux2xBits8_inst0$coreir_commonlib_mux2x8_inst0$_join_out),
		.in1(Mux2xBits8_inst1_I1_in),
		.sel(magma_Bits_8_eq_inst35_out),
		.out(Mux2xBits8_inst1$coreir_commonlib_mux2x8_inst0$_join_out)
	);
	coreir_mux #(.width(8)) Mux2xBits8_inst10$coreir_commonlib_mux2x8_inst0$_join(
		.in0(Mux2xBits8_inst9$coreir_commonlib_mux2x8_inst0$_join_out),
		.in1(Mux2xBits8_inst10_I1_in),
		.sel(magma_Bits_8_eq_inst22_out),
		.out(Mux2xBits8_inst10$coreir_commonlib_mux2x8_inst0$_join_out)
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst10_I1(
		.in(Mux2xBits8_inst10_I1_in),
		.out(a[14:7])
	);
	coreir_mux #(.width(8)) Mux2xBits8_inst11$coreir_commonlib_mux2x8_inst0$_join(
		.in0(Mux2xBits8_inst10$coreir_commonlib_mux2x8_inst0$_join_out),
		.in1(Mux2xBits8_inst11_I1_in),
		.sel(magma_Bits_8_eq_inst21_out),
		.out(Mux2xBits8_inst11$coreir_commonlib_mux2x8_inst0$_join_out)
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst11_I1(
		.in(Mux2xBits8_inst11_I1_in),
		.out(a[14:7])
	);
	coreir_mux #(.width(8)) Mux2xBits8_inst12$coreir_commonlib_mux2x8_inst0$_join(
		.in0(Mux2xBits8_inst11$coreir_commonlib_mux2x8_inst0$_join_out),
		.in1(Mux2xBits8_inst12_I1_in),
		.sel(magma_Bits_8_eq_inst20_out),
		.out(Mux2xBits8_inst12$coreir_commonlib_mux2x8_inst0$_join_out)
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst12_I1(
		.in(Mux2xBits8_inst12_I1_in),
		.out(a[14:7])
	);
	coreir_mux #(.width(8)) Mux2xBits8_inst13$coreir_commonlib_mux2x8_inst0$_join(
		.in0(Mux2xBits8_inst12$coreir_commonlib_mux2x8_inst0$_join_out),
		.in1(Mux2xBits8_inst13_I1_in),
		.sel(magma_Bits_8_eq_inst19_out),
		.out(Mux2xBits8_inst13$coreir_commonlib_mux2x8_inst0$_join_out)
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst13_I1(
		.in(Mux2xBits8_inst13_I1_in),
		.out(a[14:7])
	);
	coreir_mux #(.width(8)) Mux2xBits8_inst14$coreir_commonlib_mux2x8_inst0$_join(
		.in0(Mux2xBits8_inst13$coreir_commonlib_mux2x8_inst0$_join_out),
		.in1(Mux2xBits8_inst14_I1_in),
		.sel(magma_Bits_8_eq_inst18_out),
		.out(Mux2xBits8_inst14$coreir_commonlib_mux2x8_inst0$_join_out)
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst14_I1(
		.in(Mux2xBits8_inst14_I1_in),
		.out(a[14:7])
	);
	coreir_mux #(.width(8)) Mux2xBits8_inst15$coreir_commonlib_mux2x8_inst0$_join(
		.in0(Mux2xBits8_inst14$coreir_commonlib_mux2x8_inst0$_join_out),
		.in1(Mux2xBits8_inst15_I1_in),
		.sel(magma_Bits_8_eq_inst17_out),
		.out(Mux2xBits8_inst15$coreir_commonlib_mux2x8_inst0$_join_out)
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst15_I1(
		.in(Mux2xBits8_inst15_I1_in),
		.out(a[14:7])
	);
	coreir_mux #(.width(8)) Mux2xBits8_inst16$coreir_commonlib_mux2x8_inst0$_join(
		.in0(Mux2xBits8_inst15$coreir_commonlib_mux2x8_inst0$_join_out),
		.in1(Mux2xBits8_inst16_I1_in),
		.sel(magma_Bits_8_eq_inst16_out),
		.out(Mux2xBits8_inst16$coreir_commonlib_mux2x8_inst0$_join_out)
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst16_I1(
		.in(Mux2xBits8_inst16_I1_in),
		.out(a[14:7])
	);
	coreir_mux #(.width(8)) Mux2xBits8_inst17$coreir_commonlib_mux2x8_inst0$_join(
		.in0(Mux2xBits8_inst16$coreir_commonlib_mux2x8_inst0$_join_out),
		.in1(Mux2xBits8_inst17_I1_in),
		.sel(magma_Bits_8_eq_inst15_out),
		.out(Mux2xBits8_inst17$coreir_commonlib_mux2x8_inst0$_join_out)
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst17_I1(
		.in(Mux2xBits8_inst17_I1_in),
		.out(a[14:7])
	);
	coreir_mux #(.width(8)) Mux2xBits8_inst18$coreir_commonlib_mux2x8_inst0$_join(
		.in0(Mux2xBits8_inst17$coreir_commonlib_mux2x8_inst0$_join_out),
		.in1(Mux2xBits8_inst18_I1_in),
		.sel(magma_Bits_8_eq_inst14_out),
		.out(Mux2xBits8_inst18$coreir_commonlib_mux2x8_inst0$_join_out)
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst18_I1(
		.in(Mux2xBits8_inst18_I1_in),
		.out(a[14:7])
	);
	coreir_mux #(.width(8)) Mux2xBits8_inst19$coreir_commonlib_mux2x8_inst0$_join(
		.in0(Mux2xBits8_inst18$coreir_commonlib_mux2x8_inst0$_join_out),
		.in1(Mux2xBits8_inst19_I1_in),
		.sel(magma_Bits_8_eq_inst13_out),
		.out(Mux2xBits8_inst19$coreir_commonlib_mux2x8_inst0$_join_out)
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst19_I1(
		.in(Mux2xBits8_inst19_I1_in),
		.out(a[14:7])
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst1_I1(
		.in(Mux2xBits8_inst1_I1_in),
		.out(a[14:7])
	);
	coreir_mux #(.width(8)) Mux2xBits8_inst2$coreir_commonlib_mux2x8_inst0$_join(
		.in0(Mux2xBits8_inst1$coreir_commonlib_mux2x8_inst0$_join_out),
		.in1(Mux2xBits8_inst2_I1_in),
		.sel(magma_Bits_8_eq_inst34_out),
		.out(Mux2xBits8_inst2$coreir_commonlib_mux2x8_inst0$_join_out)
	);
	coreir_mux #(.width(8)) Mux2xBits8_inst20$coreir_commonlib_mux2x8_inst0$_join(
		.in0(Mux2xBits8_inst19$coreir_commonlib_mux2x8_inst0$_join_out),
		.in1(Mux2xBits8_inst20_I1_in),
		.sel(magma_Bit_or_inst4_out),
		.out(Mux2xBits8_inst20$coreir_commonlib_mux2x8_inst0$_join_out)
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst20_I1(
		.in(Mux2xBits8_inst20_I1_in),
		.out(a[14:7])
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst2_I1(
		.in(Mux2xBits8_inst2_I1_in),
		.out(a[14:7])
	);
	coreir_mux #(.width(8)) Mux2xBits8_inst3$coreir_commonlib_mux2x8_inst0$_join(
		.in0(Mux2xBits8_inst2$coreir_commonlib_mux2x8_inst0$_join_out),
		.in1(Mux2xBits8_inst3_I1_in),
		.sel(magma_Bits_8_eq_inst33_out),
		.out(Mux2xBits8_inst3$coreir_commonlib_mux2x8_inst0$_join_out)
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst3_I1(
		.in(Mux2xBits8_inst3_I1_in),
		.out(a[14:7])
	);
	coreir_mux #(.width(8)) Mux2xBits8_inst4$coreir_commonlib_mux2x8_inst0$_join(
		.in0(Mux2xBits8_inst3$coreir_commonlib_mux2x8_inst0$_join_out),
		.in1(Mux2xBits8_inst4_I1_in),
		.sel(magma_Bits_8_eq_inst32_out),
		.out(Mux2xBits8_inst4$coreir_commonlib_mux2x8_inst0$_join_out)
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst4_I1(
		.in(Mux2xBits8_inst4_I1_in),
		.out(a[14:7])
	);
	coreir_mux #(.width(8)) Mux2xBits8_inst5$coreir_commonlib_mux2x8_inst0$_join(
		.in0(Mux2xBits8_inst4$coreir_commonlib_mux2x8_inst0$_join_out),
		.in1(Mux2xBits8_inst5_I1_in),
		.sel(magma_Bits_8_eq_inst31_out),
		.out(Mux2xBits8_inst5$coreir_commonlib_mux2x8_inst0$_join_out)
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst5_I1(
		.in(Mux2xBits8_inst5_I1_in),
		.out(a[14:7])
	);
	coreir_mux #(.width(8)) Mux2xBits8_inst6$coreir_commonlib_mux2x8_inst0$_join(
		.in0(Mux2xBits8_inst5$coreir_commonlib_mux2x8_inst0$_join_out),
		.in1(Mux2xBits8_inst6_I1_in),
		.sel(magma_Bits_8_eq_inst30_out),
		.out(Mux2xBits8_inst6$coreir_commonlib_mux2x8_inst0$_join_out)
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst6_I1(
		.in(Mux2xBits8_inst6_I1_in),
		.out(a[14:7])
	);
	coreir_mux #(.width(8)) Mux2xBits8_inst7$coreir_commonlib_mux2x8_inst0$_join(
		.in0(Mux2xBits8_inst6$coreir_commonlib_mux2x8_inst0$_join_out),
		.in1(Mux2xBits8_inst7_I1_in),
		.sel(magma_Bit_or_inst7_out),
		.out(Mux2xBits8_inst7$coreir_commonlib_mux2x8_inst0$_join_out)
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst7_I1(
		.in(Mux2xBits8_inst7_I1_in),
		.out(a[14:7])
	);
	coreir_mux #(.width(8)) Mux2xBits8_inst8$coreir_commonlib_mux2x8_inst0$_join(
		.in0(Mux2xBits8_inst7$coreir_commonlib_mux2x8_inst0$_join_out),
		.in1(Mux2xBits8_inst8_I1_in),
		.sel(magma_Bits_8_eq_inst24_out),
		.out(Mux2xBits8_inst8$coreir_commonlib_mux2x8_inst0$_join_out)
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst8_I1(
		.in(Mux2xBits8_inst8_I1_in),
		.out(a[14:7])
	);
	coreir_mux #(.width(8)) Mux2xBits8_inst9$coreir_commonlib_mux2x8_inst0$_join(
		.in0(Mux2xBits8_inst8$coreir_commonlib_mux2x8_inst0$_join_out),
		.in1(Mux2xBits8_inst9_I1_in),
		.sel(magma_Bits_8_eq_inst23_out),
		.out(Mux2xBits8_inst9$coreir_commonlib_mux2x8_inst0$_join_out)
	);
	mantle_wire__typeBitIn8 Mux2xBits8_inst9_I1(
		.in(Mux2xBits8_inst9_I1_in),
		.out(a[14:7])
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst0$coreir_commonlib_mux2x16_inst0$_join(
		.in0(const_65409_16_out),
		.in1(const_0_16_out),
		.sel(magma_Bit_not_inst0_out),
		.out(Mux2xSInt16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst1$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst0$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_1_16_out),
		.sel(magma_Bit_not_inst1_out),
		.out(Mux2xSInt16_inst1$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst10$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst9$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_2_16_out),
		.sel(magma_Bit_not_inst11_out),
		.out(Mux2xSInt16_inst10$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst11$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst10$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_3_16_out),
		.sel(magma_Bit_not_inst12_out),
		.out(Mux2xSInt16_inst11$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst12$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst11$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_4_16_out),
		.sel(magma_Bit_not_inst13_out),
		.out(Mux2xSInt16_inst12$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst13$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst12$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_5_16_out),
		.sel(magma_Bit_not_inst14_out),
		.out(Mux2xSInt16_inst13$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst14$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst13$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_6_16_out),
		.sel(magma_Bit_not_inst15_out),
		.out(Mux2xSInt16_inst14$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst15$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst14$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_7_16_out),
		.sel(magma_Bit_not_inst16_out),
		.out(Mux2xSInt16_inst15$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst16$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst15$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_8_16_out),
		.sel(magma_Bit_not_inst17_out),
		.out(Mux2xSInt16_inst16$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst17$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst16$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_9_16_out),
		.sel(magma_Bit_not_inst18_out),
		.out(Mux2xSInt16_inst17$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst18$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst17$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_10_16_out),
		.sel(magma_Bit_not_inst19_out),
		.out(Mux2xSInt16_inst18$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst19$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst18$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_11_16_out),
		.sel(magma_Bit_not_inst20_out),
		.out(Mux2xSInt16_inst19$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst2$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst1$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_2_16_out),
		.sel(magma_Bit_not_inst2_out),
		.out(Mux2xSInt16_inst2$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst20$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst19$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_12_16_out),
		.sel(magma_Bit_not_inst21_out),
		.out(Mux2xSInt16_inst20$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst21$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst20$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_13_16_out),
		.sel(magma_Bit_not_inst22_out),
		.out(Mux2xSInt16_inst21$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst22$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst21$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_14_16_out),
		.sel(magma_Bit_not_inst23_out),
		.out(Mux2xSInt16_inst22$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst23$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst22$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_15_16_out),
		.sel(magma_Bit_not_inst24_out),
		.out(Mux2xSInt16_inst23$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst24$coreir_commonlib_mux2x16_inst0$_join(
		.in0(const_32512_16_out),
		.in1(const_127_16_out),
		.sel(magma_Bits_8_eq_inst2_out),
		.out(Mux2xSInt16_inst24$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst25$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xSInt16_inst25_I1_in),
		.sel(magma_Bits_8_eq_inst2_out),
		.out(Mux2xSInt16_inst25$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	wire [15:0] Mux2xSInt16_inst25_I1_out;
	assign Mux2xSInt16_inst25_I1_out = {Mux2xSInt9_inst0_O_out[7], Mux2xSInt9_inst0_O_out[7], Mux2xSInt9_inst0_O_out[7], Mux2xSInt9_inst0_O_out[7], Mux2xSInt9_inst0_O_out[7], Mux2xSInt9_inst0_O_out[7], Mux2xSInt9_inst0_O_out[7], Mux2xSInt9_inst0_O_out[7], Mux2xSInt9_inst0_O_out[7:0]};
	mantle_wire__typeBitIn16 Mux2xSInt16_inst25_I1(
		.in(Mux2xSInt16_inst25_I1_in),
		.out(Mux2xSInt16_inst25_I1_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst26$coreir_commonlib_mux2x16_inst0$_join(
		.in0(magma_SInt_16_sub_inst1_out),
		.in1(magma_SInt_16_sub_inst0_out),
		.sel(magma_Bits_8_eq_inst2_out),
		.out(Mux2xSInt16_inst26$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst27$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst23$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xSInt16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst2_out),
		.out(Mux2xSInt16_inst27$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst28$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst28_I0_in),
		.in1(magma_SInt_16_neg_inst2_out),
		.sel(magma_Bits_16_eq_inst0_out),
		.out(Mux2xSInt16_inst28$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	mantle_wire__typeBitIn16 Mux2xSInt16_inst28_I0(
		.in(Mux2xSInt16_inst28_I0_in),
		.out(magma_Bits_23_lshr_inst0_out[15:0])
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst29$coreir_commonlib_mux2x16_inst0$_join(
		.in0(magma_Bits_16_and_inst13_out),
		.in1(magma_SInt_16_neg_inst3_out),
		.sel(magma_Bits_16_eq_inst1_out),
		.out(Mux2xSInt16_inst29$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst3$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst2$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_3_16_out),
		.sel(magma_Bit_not_inst3_out),
		.out(Mux2xSInt16_inst3$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst30$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst29$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xSInt16_inst28$coreir_commonlib_mux2x16_inst0$_join_out),
		.sel(magma_Bits_8_eq_inst35_out),
		.out(Mux2xSInt16_inst30$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst4$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst3$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_4_16_out),
		.sel(magma_Bit_not_inst4_out),
		.out(Mux2xSInt16_inst4$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst5$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst4$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_5_16_out),
		.sel(magma_Bit_not_inst5_out),
		.out(Mux2xSInt16_inst5$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst6$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst5$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_6_16_out),
		.sel(magma_Bit_not_inst6_out),
		.out(Mux2xSInt16_inst6$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst7$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst6$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_7_16_out),
		.sel(magma_Bit_not_inst7_out),
		.out(Mux2xSInt16_inst7$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst8$coreir_commonlib_mux2x16_inst0$_join(
		.in0(const_65409_16_out),
		.in1(const_0_16_out),
		.sel(magma_Bit_not_inst9_out),
		.out(Mux2xSInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(16)) Mux2xSInt16_inst9$coreir_commonlib_mux2x16_inst0$_join(
		.in0(Mux2xSInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_1_16_out),
		.sel(magma_Bit_not_inst10_out),
		.out(Mux2xSInt16_inst9$coreir_commonlib_mux2x16_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst0$coreir_commonlib_mux2x9_inst0$_join(
		.in0(magma_SInt_9_sub_inst0_out),
		.in1(magma_SInt_9_neg_inst0_out),
		.sel(magma_SInt_9_slt_inst0_out),
		.out(Mux2xSInt9_inst0$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	mantle_wire__typeBit9 Mux2xSInt9_inst0_O(
		.in(Mux2xSInt9_inst0$coreir_commonlib_mux2x9_inst0$_join_out),
		.out(Mux2xSInt9_inst0_O_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst1$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst1_I0_in),
		.in1(Mux2xSInt9_inst1_I1_in),
		.sel(magma_Bits_8_eq_inst36_out),
		.out(Mux2xSInt9_inst1$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst10$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst8$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(magma_SInt_9_sub_inst0_out),
		.sel(magma_Bits_8_eq_inst32_out),
		.out(Mux2xSInt9_inst10$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst11$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst9$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(Mux2xSInt9_inst11_I1_in),
		.sel(magma_Bits_8_eq_inst31_out),
		.out(Mux2xSInt9_inst11$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	wire [8:0] Mux2xSInt9_inst11_I1_out;
	assign Mux2xSInt9_inst11_I1_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst11_I1(
		.in(Mux2xSInt9_inst11_I1_in),
		.out(Mux2xSInt9_inst11_I1_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst12$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst10$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(magma_SInt_9_sub_inst0_out),
		.sel(magma_Bits_8_eq_inst31_out),
		.out(Mux2xSInt9_inst12$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst13$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst11$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(Mux2xSInt9_inst13_I1_in),
		.sel(magma_Bits_8_eq_inst30_out),
		.out(Mux2xSInt9_inst13$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	wire [8:0] Mux2xSInt9_inst13_I1_out;
	assign Mux2xSInt9_inst13_I1_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst13_I1(
		.in(Mux2xSInt9_inst13_I1_in),
		.out(Mux2xSInt9_inst13_I1_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst14$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst12$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(magma_SInt_9_sub_inst0_out),
		.sel(magma_Bits_8_eq_inst30_out),
		.out(Mux2xSInt9_inst14$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst15$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst13$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(Mux2xSInt9_inst15_I1_in),
		.sel(magma_Bit_or_inst7_out),
		.out(Mux2xSInt9_inst15$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	wire [8:0] Mux2xSInt9_inst15_I1_out;
	assign Mux2xSInt9_inst15_I1_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst15_I1(
		.in(Mux2xSInt9_inst15_I1_in),
		.out(Mux2xSInt9_inst15_I1_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst16$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst14$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(magma_SInt_9_sub_inst0_out),
		.sel(magma_Bit_or_inst7_out),
		.out(Mux2xSInt9_inst16$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst17$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst15$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(Mux2xSInt9_inst17_I1_in),
		.sel(magma_Bits_8_eq_inst24_out),
		.out(Mux2xSInt9_inst17$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	wire [8:0] Mux2xSInt9_inst17_I1_out;
	assign Mux2xSInt9_inst17_I1_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst17_I1(
		.in(Mux2xSInt9_inst17_I1_in),
		.out(Mux2xSInt9_inst17_I1_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst18$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst16$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(magma_SInt_9_sub_inst0_out),
		.sel(magma_Bits_8_eq_inst24_out),
		.out(Mux2xSInt9_inst18$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst19$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst17$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(Mux2xSInt9_inst19_I1_in),
		.sel(magma_Bits_8_eq_inst23_out),
		.out(Mux2xSInt9_inst19$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	wire [8:0] Mux2xSInt9_inst19_I1_out;
	assign Mux2xSInt9_inst19_I1_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst19_I1(
		.in(Mux2xSInt9_inst19_I1_in),
		.out(Mux2xSInt9_inst19_I1_out)
	);
	wire [8:0] Mux2xSInt9_inst1_I0_out;
	assign Mux2xSInt9_inst1_I0_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst1_I0(
		.in(Mux2xSInt9_inst1_I0_in),
		.out(Mux2xSInt9_inst1_I0_out)
	);
	wire [8:0] Mux2xSInt9_inst1_I1_out;
	assign Mux2xSInt9_inst1_I1_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst1_I1(
		.in(Mux2xSInt9_inst1_I1_in),
		.out(Mux2xSInt9_inst1_I1_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst2$coreir_commonlib_mux2x9_inst0$_join(
		.in0(magma_SInt_9_sub_inst0_out),
		.in1(magma_SInt_9_sub_inst2_out),
		.sel(magma_Bits_8_eq_inst36_out),
		.out(Mux2xSInt9_inst2$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst20$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst18$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(magma_SInt_9_sub_inst0_out),
		.sel(magma_Bits_8_eq_inst23_out),
		.out(Mux2xSInt9_inst20$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst21$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst19$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(Mux2xSInt9_inst21_I1_in),
		.sel(magma_Bits_8_eq_inst22_out),
		.out(Mux2xSInt9_inst21$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	wire [8:0] Mux2xSInt9_inst21_I1_out;
	assign Mux2xSInt9_inst21_I1_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst21_I1(
		.in(Mux2xSInt9_inst21_I1_in),
		.out(Mux2xSInt9_inst21_I1_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst22$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst20$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(magma_SInt_9_sub_inst0_out),
		.sel(magma_Bits_8_eq_inst22_out),
		.out(Mux2xSInt9_inst22$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst23$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst21$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(Mux2xSInt9_inst23_I1_in),
		.sel(magma_Bits_8_eq_inst21_out),
		.out(Mux2xSInt9_inst23$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	wire [8:0] Mux2xSInt9_inst23_I1_out;
	assign Mux2xSInt9_inst23_I1_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst23_I1(
		.in(Mux2xSInt9_inst23_I1_in),
		.out(Mux2xSInt9_inst23_I1_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst24$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst22$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(magma_SInt_9_sub_inst0_out),
		.sel(magma_Bits_8_eq_inst21_out),
		.out(Mux2xSInt9_inst24$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst25$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst23$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(Mux2xSInt9_inst25_I1_in),
		.sel(magma_Bits_8_eq_inst20_out),
		.out(Mux2xSInt9_inst25$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	wire [8:0] Mux2xSInt9_inst25_I1_out;
	assign Mux2xSInt9_inst25_I1_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst25_I1(
		.in(Mux2xSInt9_inst25_I1_in),
		.out(Mux2xSInt9_inst25_I1_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst26$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst24$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(magma_SInt_9_sub_inst0_out),
		.sel(magma_Bits_8_eq_inst20_out),
		.out(Mux2xSInt9_inst26$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst27$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst25$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(Mux2xSInt9_inst27_I1_in),
		.sel(magma_Bits_8_eq_inst19_out),
		.out(Mux2xSInt9_inst27$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	wire [8:0] Mux2xSInt9_inst27_I1_out;
	assign Mux2xSInt9_inst27_I1_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst27_I1(
		.in(Mux2xSInt9_inst27_I1_in),
		.out(Mux2xSInt9_inst27_I1_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst28$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst26$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(magma_SInt_9_sub_inst0_out),
		.sel(magma_Bits_8_eq_inst19_out),
		.out(Mux2xSInt9_inst28$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst29$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst27$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(Mux2xSInt9_inst29_I1_in),
		.sel(magma_Bits_8_eq_inst18_out),
		.out(Mux2xSInt9_inst29$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	wire [8:0] Mux2xSInt9_inst29_I1_out;
	assign Mux2xSInt9_inst29_I1_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst29_I1(
		.in(Mux2xSInt9_inst29_I1_in),
		.out(Mux2xSInt9_inst29_I1_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst3$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst1$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(Mux2xSInt9_inst3_I1_in),
		.sel(magma_Bits_8_eq_inst35_out),
		.out(Mux2xSInt9_inst3$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst30$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst28$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(magma_SInt_9_sub_inst0_out),
		.sel(magma_Bits_8_eq_inst18_out),
		.out(Mux2xSInt9_inst30$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst31$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst29$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(Mux2xSInt9_inst31_I1_in),
		.sel(magma_Bits_8_eq_inst17_out),
		.out(Mux2xSInt9_inst31$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	wire [8:0] Mux2xSInt9_inst31_I1_out;
	assign Mux2xSInt9_inst31_I1_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst31_I1(
		.in(Mux2xSInt9_inst31_I1_in),
		.out(Mux2xSInt9_inst31_I1_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst32$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst30$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(magma_SInt_9_sub_inst0_out),
		.sel(magma_Bits_8_eq_inst17_out),
		.out(Mux2xSInt9_inst32$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst33$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst31$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(Mux2xSInt9_inst33_I1_in),
		.sel(magma_Bits_8_eq_inst16_out),
		.out(Mux2xSInt9_inst33$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	wire [8:0] Mux2xSInt9_inst33_I1_out;
	assign Mux2xSInt9_inst33_I1_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst33_I1(
		.in(Mux2xSInt9_inst33_I1_in),
		.out(Mux2xSInt9_inst33_I1_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst34$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst32$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(magma_SInt_9_sub_inst0_out),
		.sel(magma_Bits_8_eq_inst16_out),
		.out(Mux2xSInt9_inst34$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst35$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst33$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(Mux2xSInt9_inst35_I1_in),
		.sel(magma_Bits_8_eq_inst15_out),
		.out(Mux2xSInt9_inst35$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	wire [8:0] Mux2xSInt9_inst35_I1_out;
	assign Mux2xSInt9_inst35_I1_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst35_I1(
		.in(Mux2xSInt9_inst35_I1_in),
		.out(Mux2xSInt9_inst35_I1_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst36$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst34$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(magma_SInt_9_sub_inst0_out),
		.sel(magma_Bits_8_eq_inst15_out),
		.out(Mux2xSInt9_inst36$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst37$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst35$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(Mux2xSInt9_inst37_I1_in),
		.sel(magma_Bits_8_eq_inst14_out),
		.out(Mux2xSInt9_inst37$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	wire [8:0] Mux2xSInt9_inst37_I1_out;
	assign Mux2xSInt9_inst37_I1_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst37_I1(
		.in(Mux2xSInt9_inst37_I1_in),
		.out(Mux2xSInt9_inst37_I1_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst38$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst36$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(magma_SInt_9_sub_inst0_out),
		.sel(magma_Bits_8_eq_inst14_out),
		.out(Mux2xSInt9_inst38$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst39$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst37$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(Mux2xSInt9_inst39_I1_in),
		.sel(magma_Bits_8_eq_inst13_out),
		.out(Mux2xSInt9_inst39$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	wire [8:0] Mux2xSInt9_inst39_I1_out;
	assign Mux2xSInt9_inst39_I1_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst39_I1(
		.in(Mux2xSInt9_inst39_I1_in),
		.out(Mux2xSInt9_inst39_I1_out)
	);
	wire [8:0] Mux2xSInt9_inst3_I1_out;
	assign Mux2xSInt9_inst3_I1_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst3_I1(
		.in(Mux2xSInt9_inst3_I1_in),
		.out(Mux2xSInt9_inst3_I1_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst4$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst2$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(magma_SInt_9_sub_inst1_out),
		.sel(magma_Bits_8_eq_inst35_out),
		.out(Mux2xSInt9_inst4$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst40$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst38$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(magma_SInt_9_sub_inst0_out),
		.sel(magma_Bits_8_eq_inst13_out),
		.out(Mux2xSInt9_inst40$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst41$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst39$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(Mux2xSInt9_inst41_I1_in),
		.sel(magma_Bit_or_inst4_out),
		.out(Mux2xSInt9_inst41$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	wire [8:0] Mux2xSInt9_inst41_I1_out;
	assign Mux2xSInt9_inst41_I1_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst41_I1(
		.in(Mux2xSInt9_inst41_I1_in),
		.out(Mux2xSInt9_inst41_I1_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst42$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst40$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(magma_SInt_9_sub_inst0_out),
		.sel(magma_Bit_or_inst4_out),
		.out(Mux2xSInt9_inst42$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst5$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst3$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(Mux2xSInt9_inst5_I1_in),
		.sel(magma_Bits_8_eq_inst34_out),
		.out(Mux2xSInt9_inst5$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	wire [8:0] Mux2xSInt9_inst5_I1_out;
	assign Mux2xSInt9_inst5_I1_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst5_I1(
		.in(Mux2xSInt9_inst5_I1_in),
		.out(Mux2xSInt9_inst5_I1_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst6$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst4$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(magma_SInt_9_sub_inst0_out),
		.sel(magma_Bits_8_eq_inst34_out),
		.out(Mux2xSInt9_inst6$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst7$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst5$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(Mux2xSInt9_inst7_I1_in),
		.sel(magma_Bits_8_eq_inst33_out),
		.out(Mux2xSInt9_inst7$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	wire [8:0] Mux2xSInt9_inst7_I1_out;
	assign Mux2xSInt9_inst7_I1_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst7_I1(
		.in(Mux2xSInt9_inst7_I1_in),
		.out(Mux2xSInt9_inst7_I1_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst8$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst6$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(magma_SInt_9_sub_inst0_out),
		.sel(magma_Bits_8_eq_inst33_out),
		.out(Mux2xSInt9_inst8$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	coreir_mux #(.width(9)) Mux2xSInt9_inst9$coreir_commonlib_mux2x9_inst0$_join(
		.in0(Mux2xSInt9_inst7$coreir_commonlib_mux2x9_inst0$_join_out),
		.in1(Mux2xSInt9_inst9_I1_in),
		.sel(magma_Bits_8_eq_inst32_out),
		.out(Mux2xSInt9_inst9$coreir_commonlib_mux2x9_inst0$_join_out)
	);
	wire [8:0] Mux2xSInt9_inst9_I1_out;
	assign Mux2xSInt9_inst9_I1_out = {bit_const_0_None_out, a[14:7]};
	mantle_wire__typeBitIn9 Mux2xSInt9_inst9_I1(
		.in(Mux2xSInt9_inst9_I1_in),
		.out(Mux2xSInt9_inst9_I1_out)
	);
	coreir_mux #(.width(32)) Mux2xUInt32_inst0$coreir_commonlib_mux2x32_inst0$_join(
		.in0(Mux2xUInt32_inst0_I0_in),
		.in1(Mux2xUInt32_inst0_I1_in),
		.sel(magma_Bits_1_eq_inst0_out),
		.out(Mux2xUInt32_inst0$coreir_commonlib_mux2x32_inst0$_join_out)
	);
	wire [31:0] Mux2xUInt32_inst0_I0_out;
	assign Mux2xUInt32_inst0_I0_out = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, a[15:0]};
	mantle_wire__typeBitIn32 Mux2xUInt32_inst0_I0(
		.in(Mux2xUInt32_inst0_I0_in),
		.out(Mux2xUInt32_inst0_I0_out)
	);
	wire [31:0] Mux2xUInt32_inst0_I1_out;
	assign Mux2xUInt32_inst0_I1_out = {a[15], a[15], a[15], a[15], a[15], a[15], a[15], a[15], a[15], a[15], a[15], a[15], a[15], a[15], a[15], a[15], a[15:0]};
	mantle_wire__typeBitIn32 Mux2xUInt32_inst0_I1(
		.in(Mux2xUInt32_inst0_I1_in),
		.out(Mux2xUInt32_inst0_I1_out)
	);
	coreir_mux #(.width(32)) Mux2xUInt32_inst1$coreir_commonlib_mux2x32_inst0$_join(
		.in0(Mux2xUInt32_inst1_I0_in),
		.in1(Mux2xUInt32_inst1_I1_in),
		.sel(magma_Bits_1_eq_inst0_out),
		.out(Mux2xUInt32_inst1$coreir_commonlib_mux2x32_inst0$_join_out)
	);
	wire [31:0] Mux2xUInt32_inst1_I0_out;
	assign Mux2xUInt32_inst1_I0_out = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, b[15:0]};
	mantle_wire__typeBitIn32 Mux2xUInt32_inst1_I0(
		.in(Mux2xUInt32_inst1_I0_in),
		.out(Mux2xUInt32_inst1_I0_out)
	);
	wire [31:0] Mux2xUInt32_inst1_I1_out;
	assign Mux2xUInt32_inst1_I1_out = {b[15], b[15], b[15], b[15], b[15], b[15], b[15], b[15], b[15], b[15], b[15], b[15], b[15], b[15], b[15], b[15], b[15:0]};
	mantle_wire__typeBitIn32 Mux2xUInt32_inst1_I1(
		.in(Mux2xUInt32_inst1_I1_in),
		.out(Mux2xUInt32_inst1_I1_out)
	);
	corebit_const #(.value(1'b0)) bit_const_0_None(.out(bit_const_0_None_out));
	corebit_const #(.value(1'b1)) bit_const_1_None(.out(bit_const_1_None_out));
	coreir_const #(
		.value(16'h0000),
		.width(16)
	) const_0_16(.out(const_0_16_out));
	coreir_const #(
		.value(23'h000000),
		.width(23)
	) const_0_23(.out(const_0_23_out));
	coreir_const #(
		.value(7'h00),
		.width(7)
	) const_0_7(.out(const_0_7_out));
	coreir_const #(
		.value(8'h00),
		.width(8)
	) const_0_8(.out(const_0_8_out));
	coreir_const #(
		.value(9'h000),
		.width(9)
	) const_0_9(.out(const_0_9_out));
	coreir_const #(
		.value(16'h000a),
		.width(16)
	) const_10_16(.out(const_10_16_out));
	coreir_const #(
		.value(16'h000b),
		.width(16)
	) const_11_16(.out(const_11_16_out));
	coreir_const #(
		.value(8'h0b),
		.width(8)
	) const_11_8(.out(const_11_8_out));
	coreir_const #(
		.value(16'h007f),
		.width(16)
	) const_127_16(.out(const_127_16_out));
	coreir_const #(
		.value(8'h7f),
		.width(8)
	) const_127_8(.out(const_127_8_out));
	coreir_const #(
		.value(9'h07f),
		.width(9)
	) const_127_9(.out(const_127_9_out));
	coreir_const #(
		.value(16'h0080),
		.width(16)
	) const_128_16(.out(const_128_16_out));
	coreir_const #(
		.value(16'h000c),
		.width(16)
	) const_12_16(.out(const_12_16_out));
	coreir_const #(
		.value(8'h0c),
		.width(8)
	) const_12_8(.out(const_12_8_out));
	coreir_const #(
		.value(16'h000d),
		.width(16)
	) const_13_16(.out(const_13_16_out));
	coreir_const #(
		.value(8'h0d),
		.width(8)
	) const_13_8(.out(const_13_8_out));
	coreir_const #(
		.value(8'h8e),
		.width(8)
	) const_142_8(.out(const_142_8_out));
	coreir_const #(
		.value(8'h92),
		.width(8)
	) const_146_8(.out(const_146_8_out));
	coreir_const #(
		.value(8'h93),
		.width(8)
	) const_147_8(.out(const_147_8_out));
	coreir_const #(
		.value(8'h94),
		.width(8)
	) const_148_8(.out(const_148_8_out));
	coreir_const #(
		.value(8'h95),
		.width(8)
	) const_149_8(.out(const_149_8_out));
	coreir_const #(
		.value(16'h000e),
		.width(16)
	) const_14_16(.out(const_14_16_out));
	coreir_const #(
		.value(8'h96),
		.width(8)
	) const_150_8(.out(const_150_8_out));
	coreir_const #(
		.value(8'h97),
		.width(8)
	) const_151_8(.out(const_151_8_out));
	coreir_const #(
		.value(8'h98),
		.width(8)
	) const_152_8(.out(const_152_8_out));
	coreir_const #(
		.value(16'h000f),
		.width(16)
	) const_15_16(.out(const_15_16_out));
	coreir_const #(
		.value(8'h0f),
		.width(8)
	) const_15_8(.out(const_15_8_out));
	coreir_const #(
		.value(8'h11),
		.width(8)
	) const_17_8(.out(const_17_8_out));
	coreir_const #(
		.value(8'h12),
		.width(8)
	) const_18_8(.out(const_18_8_out));
	coreir_const #(
		.value(8'h13),
		.width(8)
	) const_19_8(.out(const_19_8_out));
	coreir_const #(
		.value(1'h1),
		.width(1)
	) const_1_1(.out(const_1_1_out));
	coreir_const #(
		.value(16'h0001),
		.width(16)
	) const_1_16(.out(const_1_16_out));
	coreir_const #(
		.value(8'h01),
		.width(8)
	) const_1_8(.out(const_1_8_out));
	coreir_const #(
		.value(8'h14),
		.width(8)
	) const_20_8(.out(const_20_8_out));
	coreir_const #(
		.value(8'h16),
		.width(8)
	) const_22_8(.out(const_22_8_out));
	coreir_const #(
		.value(8'h17),
		.width(8)
	) const_23_8(.out(const_23_8_out));
	coreir_const #(
		.value(8'h18),
		.width(8)
	) const_24_8(.out(const_24_8_out));
	coreir_const #(
		.value(8'hff),
		.width(8)
	) const_255_8(.out(const_255_8_out));
	coreir_const #(
		.value(9'h0ff),
		.width(9)
	) const_255_9(.out(const_255_9_out));
	coreir_const #(
		.value(8'h19),
		.width(8)
	) const_25_8(.out(const_25_8_out));
	coreir_const #(
		.value(16'h0002),
		.width(16)
	) const_2_16(.out(const_2_16_out));
	coreir_const #(
		.value(8'h02),
		.width(8)
	) const_2_8(.out(const_2_8_out));
	coreir_const #(
		.value(16'h7f00),
		.width(16)
	) const_32512_16(.out(const_32512_16_out));
	coreir_const #(
		.value(16'h7f80),
		.width(16)
	) const_32640_16(.out(const_32640_16_out));
	coreir_const #(
		.value(16'h8000),
		.width(16)
	) const_32768_16(.out(const_32768_16_out));
	coreir_const #(
		.value(16'h0003),
		.width(16)
	) const_3_16(.out(const_3_16_out));
	coreir_const #(
		.value(8'h03),
		.width(8)
	) const_3_8(.out(const_3_8_out));
	coreir_const #(
		.value(16'h0004),
		.width(16)
	) const_4_16(.out(const_4_16_out));
	coreir_const #(
		.value(8'h04),
		.width(8)
	) const_4_8(.out(const_4_8_out));
	coreir_const #(
		.value(16'h0005),
		.width(16)
	) const_5_16(.out(const_5_16_out));
	coreir_const #(
		.value(8'h05),
		.width(8)
	) const_5_8(.out(const_5_8_out));
	coreir_const #(
		.value(16'hff81),
		.width(16)
	) const_65409_16(.out(const_65409_16_out));
	coreir_const #(
		.value(16'h0006),
		.width(16)
	) const_6_16(.out(const_6_16_out));
	coreir_const #(
		.value(8'h06),
		.width(8)
	) const_6_8(.out(const_6_8_out));
	coreir_const #(
		.value(16'h0007),
		.width(16)
	) const_7_16(.out(const_7_16_out));
	coreir_const #(
		.value(23'h000007),
		.width(23)
	) const_7_23(.out(const_7_23_out));
	coreir_const #(
		.value(16'h0008),
		.width(16)
	) const_8_16(.out(const_8_16_out));
	coreir_const #(
		.value(8'h08),
		.width(8)
	) const_8_8(.out(const_8_8_out));
	coreir_const #(
		.value(16'h0009),
		.width(16)
	) const_9_16(.out(const_9_16_out));
	assign magma_BFloat_16_mul_inst0_out = 16'd0;
	assign magma_BFloat_16_add_inst0_out = 16'd0;
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_8_eq_inst0_out),
		.in1(magma_Bits_7_eq_inst0_out),
		.out(magma_Bit_and_inst0_out)
	);
	corebit_and magma_Bit_and_inst1(
		.in0(magma_Bits_8_eq_inst1_out),
		.in1(magma_Bits_7_eq_inst1_out),
		.out(magma_Bit_and_inst1_out)
	);
	corebit_and magma_Bit_and_inst2(
		.in0(a[15]),
		.in1(Mux2xBits16_inst7_O_out[15]),
		.out(magma_Bit_and_inst2_out)
	);
	corebit_and magma_Bit_and_inst3(
		.in0(magma_Bit_and_inst2_out),
		.in1(magma_Bit_not_inst25_out),
		.out(magma_Bit_and_inst3_out)
	);
	corebit_and magma_Bit_and_inst4(
		.in0(magma_Bit_not_inst26_out),
		.in1(magma_Bit_not_inst27_out),
		.out(magma_Bit_and_inst4_out)
	);
	corebit_and magma_Bit_and_inst5(
		.in0(magma_Bit_and_inst4_out),
		.in1(magma_UInt_17_add_inst1_out[15]),
		.out(magma_Bit_and_inst5_out)
	);
	corebit_and magma_Bit_and_inst6(
		.in0(magma_Bits_8_eq_inst41_out),
		.in1(magma_Bits_7_eq_inst2_out),
		.out(magma_Bit_and_inst6_out)
	);
	corebit_and magma_Bit_and_inst7(
		.in0(magma_Bit_and_inst0_out),
		.in1(magma_Bit_and_inst1_out),
		.out(magma_Bit_and_inst7_out)
	);
	corebit_and magma_Bit_and_inst8(
		.in0(magma_Bit_and_inst7_out),
		.in1(magma_Bit_not_inst28_out),
		.out(magma_Bit_and_inst8_out)
	);
	corebit_not magma_Bit_not_inst0(
		.in(magma_Bit_xor_inst0_out),
		.out(magma_Bit_not_inst0_out)
	);
	corebit_not magma_Bit_not_inst1(
		.in(magma_Bit_xor_inst1_out),
		.out(magma_Bit_not_inst1_out)
	);
	corebit_not magma_Bit_not_inst10(
		.in(magma_Bit_xor_inst10_out),
		.out(magma_Bit_not_inst10_out)
	);
	corebit_not magma_Bit_not_inst11(
		.in(magma_Bit_xor_inst11_out),
		.out(magma_Bit_not_inst11_out)
	);
	corebit_not magma_Bit_not_inst12(
		.in(magma_Bit_xor_inst12_out),
		.out(magma_Bit_not_inst12_out)
	);
	corebit_not magma_Bit_not_inst13(
		.in(magma_Bit_xor_inst13_out),
		.out(magma_Bit_not_inst13_out)
	);
	corebit_not magma_Bit_not_inst14(
		.in(magma_Bit_xor_inst14_out),
		.out(magma_Bit_not_inst14_out)
	);
	corebit_not magma_Bit_not_inst15(
		.in(magma_Bit_xor_inst15_out),
		.out(magma_Bit_not_inst15_out)
	);
	corebit_not magma_Bit_not_inst16(
		.in(magma_Bit_xor_inst16_out),
		.out(magma_Bit_not_inst16_out)
	);
	corebit_not magma_Bit_not_inst17(
		.in(magma_Bit_xor_inst17_out),
		.out(magma_Bit_not_inst17_out)
	);
	corebit_not magma_Bit_not_inst18(
		.in(magma_Bit_xor_inst18_out),
		.out(magma_Bit_not_inst18_out)
	);
	corebit_not magma_Bit_not_inst19(
		.in(magma_Bit_xor_inst19_out),
		.out(magma_Bit_not_inst19_out)
	);
	corebit_not magma_Bit_not_inst2(
		.in(magma_Bit_xor_inst2_out),
		.out(magma_Bit_not_inst2_out)
	);
	corebit_not magma_Bit_not_inst20(
		.in(magma_Bit_xor_inst20_out),
		.out(magma_Bit_not_inst20_out)
	);
	corebit_not magma_Bit_not_inst21(
		.in(magma_Bit_xor_inst21_out),
		.out(magma_Bit_not_inst21_out)
	);
	corebit_not magma_Bit_not_inst22(
		.in(magma_Bit_xor_inst22_out),
		.out(magma_Bit_not_inst22_out)
	);
	corebit_not magma_Bit_not_inst23(
		.in(magma_Bit_xor_inst23_out),
		.out(magma_Bit_not_inst23_out)
	);
	corebit_not magma_Bit_not_inst24(
		.in(magma_Bit_xor_inst24_out),
		.out(magma_Bit_not_inst24_out)
	);
	corebit_not magma_Bit_not_inst25(
		.in(magma_UInt_17_add_inst1_out[15]),
		.out(magma_Bit_not_inst25_out)
	);
	corebit_not magma_Bit_not_inst26(
		.in(a[15]),
		.out(magma_Bit_not_inst26_out)
	);
	corebit_not magma_Bit_not_inst27(
		.in(Mux2xBits16_inst7_O_out[15]),
		.out(magma_Bit_not_inst27_out)
	);
	corebit_not magma_Bit_not_inst28(
		.in(magma_Bit_xor_inst25_out),
		.out(magma_Bit_not_inst28_out)
	);
	corebit_not magma_Bit_not_inst3(
		.in(magma_Bit_xor_inst3_out),
		.out(magma_Bit_not_inst3_out)
	);
	corebit_not magma_Bit_not_inst4(
		.in(magma_Bit_xor_inst4_out),
		.out(magma_Bit_not_inst4_out)
	);
	corebit_not magma_Bit_not_inst5(
		.in(magma_Bit_xor_inst5_out),
		.out(magma_Bit_not_inst5_out)
	);
	corebit_not magma_Bit_not_inst6(
		.in(magma_Bit_xor_inst6_out),
		.out(magma_Bit_not_inst6_out)
	);
	corebit_not magma_Bit_not_inst7(
		.in(magma_Bit_xor_inst7_out),
		.out(magma_Bit_not_inst7_out)
	);
	corebit_not magma_Bit_not_inst8(
		.in(magma_Bit_xor_inst8_out),
		.out(magma_Bit_not_inst8_out)
	);
	corebit_not magma_Bit_not_inst9(
		.in(magma_Bit_xor_inst9_out),
		.out(magma_Bit_not_inst9_out)
	);
	corebit_or magma_Bit_or_inst0(
		.in0(magma_Bits_8_eq_inst4_out),
		.in1(magma_Bits_8_eq_inst5_out),
		.out(magma_Bit_or_inst0_out)
	);
	corebit_or magma_Bit_or_inst1(
		.in0(magma_Bits_8_eq_inst7_out),
		.in1(magma_Bits_8_eq_inst8_out),
		.out(magma_Bit_or_inst1_out)
	);
	corebit_or magma_Bit_or_inst10(
		.in0(magma_Bit_or_inst9_out),
		.in1(magma_Bits_8_eq_inst39_out),
		.out(magma_Bit_or_inst10_out)
	);
	corebit_or magma_Bit_or_inst11(
		.in0(magma_Bit_or_inst10_out),
		.in1(magma_Bits_8_eq_inst40_out),
		.out(magma_Bit_or_inst11_out)
	);
	corebit_or magma_Bit_or_inst12(
		.in0(magma_Bits_8_eq_inst14_out),
		.in1(magma_Bits_8_eq_inst15_out),
		.out(magma_Bit_or_inst12_out)
	);
	corebit_or magma_Bit_or_inst13(
		.in0(magma_Bit_or_inst12_out),
		.in1(magma_Bits_8_eq_inst13_out),
		.out(magma_Bit_or_inst13_out)
	);
	corebit_or magma_Bit_or_inst2(
		.in0(magma_Bits_8_eq_inst9_out),
		.in1(magma_Bits_8_eq_inst10_out),
		.out(magma_Bit_or_inst2_out)
	);
	corebit_or magma_Bit_or_inst3(
		.in0(magma_Bit_or_inst2_out),
		.in1(magma_Bits_8_eq_inst11_out),
		.out(magma_Bit_or_inst3_out)
	);
	corebit_or magma_Bit_or_inst4(
		.in0(magma_Bit_or_inst3_out),
		.in1(magma_Bits_8_eq_inst12_out),
		.out(magma_Bit_or_inst4_out)
	);
	corebit_or magma_Bit_or_inst5(
		.in0(magma_Bit_and_inst3_out),
		.in1(magma_Bit_and_inst5_out),
		.out(magma_Bit_or_inst5_out)
	);
	corebit_or magma_Bit_or_inst6(
		.in0(magma_Bits_8_eq_inst25_out),
		.in1(magma_Bits_8_eq_inst26_out),
		.out(magma_Bit_or_inst6_out)
	);
	corebit_or magma_Bit_or_inst7(
		.in0(magma_Bit_or_inst6_out),
		.in1(magma_Bits_8_eq_inst27_out),
		.out(magma_Bit_or_inst7_out)
	);
	corebit_or magma_Bit_or_inst8(
		.in0(magma_Bits_8_eq_inst28_out),
		.in1(magma_Bits_8_eq_inst29_out),
		.out(magma_Bit_or_inst8_out)
	);
	corebit_or magma_Bit_or_inst9(
		.in0(magma_Bits_8_eq_inst37_out),
		.in1(magma_Bits_8_eq_inst38_out),
		.out(magma_Bit_or_inst9_out)
	);
	corebit_xor magma_Bit_xor_inst0(
		.in0(Mux2xSInt9_inst0_O_out[0]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst0_out)
	);
	corebit_xor magma_Bit_xor_inst1(
		.in0(Mux2xSInt9_inst0_O_out[1]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst1_out)
	);
	corebit_xor magma_Bit_xor_inst10(
		.in0(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out[1]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst10_out)
	);
	corebit_xor magma_Bit_xor_inst11(
		.in0(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out[2]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst11_out)
	);
	corebit_xor magma_Bit_xor_inst12(
		.in0(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out[3]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst12_out)
	);
	corebit_xor magma_Bit_xor_inst13(
		.in0(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out[4]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst13_out)
	);
	corebit_xor magma_Bit_xor_inst14(
		.in0(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out[5]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst14_out)
	);
	corebit_xor magma_Bit_xor_inst15(
		.in0(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out[6]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst15_out)
	);
	corebit_xor magma_Bit_xor_inst16(
		.in0(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out[7]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst16_out)
	);
	corebit_xor magma_Bit_xor_inst17(
		.in0(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out[8]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst17_out)
	);
	corebit_xor magma_Bit_xor_inst18(
		.in0(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out[9]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst18_out)
	);
	corebit_xor magma_Bit_xor_inst19(
		.in0(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out[10]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst19_out)
	);
	corebit_xor magma_Bit_xor_inst2(
		.in0(Mux2xSInt9_inst0_O_out[2]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst2_out)
	);
	corebit_xor magma_Bit_xor_inst20(
		.in0(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out[11]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst20_out)
	);
	corebit_xor magma_Bit_xor_inst21(
		.in0(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out[12]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst21_out)
	);
	corebit_xor magma_Bit_xor_inst22(
		.in0(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out[13]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst22_out)
	);
	corebit_xor magma_Bit_xor_inst23(
		.in0(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out[14]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst23_out)
	);
	corebit_xor magma_Bit_xor_inst24(
		.in0(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out[15]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst24_out)
	);
	corebit_xor magma_Bit_xor_inst25(
		.in0(a[15]),
		.in1(b[15]),
		.out(magma_Bit_xor_inst25_out)
	);
	corebit_xor magma_Bit_xor_inst3(
		.in0(Mux2xSInt9_inst0_O_out[3]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst3_out)
	);
	corebit_xor magma_Bit_xor_inst4(
		.in0(Mux2xSInt9_inst0_O_out[4]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst4_out)
	);
	corebit_xor magma_Bit_xor_inst5(
		.in0(Mux2xSInt9_inst0_O_out[5]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst5_out)
	);
	corebit_xor magma_Bit_xor_inst6(
		.in0(Mux2xSInt9_inst0_O_out[6]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst6_out)
	);
	corebit_xor magma_Bit_xor_inst7(
		.in0(Mux2xSInt9_inst0_O_out[7]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst7_out)
	);
	corebit_xor magma_Bit_xor_inst8(
		.in0(Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_out[15]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst8_out)
	);
	corebit_xor magma_Bit_xor_inst9(
		.in0(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out[0]),
		.in1(bit_const_1_None_out),
		.out(magma_Bit_xor_inst9_out)
	);
	coreir_and #(.width(16)) magma_Bits_16_and_inst0(
		.in0(a),
		.in1(const_32768_16_out),
		.out(magma_Bits_16_and_inst0_out)
	);
	coreir_and #(.width(16)) magma_Bits_16_and_inst1(
		.in0(magma_Bits_16_shl_inst0_out),
		.in1(const_32640_16_out),
		.out(magma_Bits_16_and_inst1_out)
	);
	coreir_and #(.width(16)) magma_Bits_16_and_inst10(
		.in0(a),
		.in1(const_127_16_out),
		.out(magma_Bits_16_and_inst10_out)
	);
	coreir_and #(.width(16)) magma_Bits_16_and_inst11(
		.in0(a),
		.in1(const_32768_16_out),
		.out(magma_Bits_16_and_inst11_out)
	);
	coreir_and #(.width(16)) magma_Bits_16_and_inst12(
		.in0(a),
		.in1(const_127_16_out),
		.out(magma_Bits_16_and_inst12_out)
	);
	coreir_and #(.width(16)) magma_Bits_16_and_inst13(
		.in0(Mux2xBits16_inst13$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_127_16_out),
		.out(magma_Bits_16_and_inst13_out)
	);
	wire [15:0] magma_Bits_16_and_inst14_in1;
	assign magma_Bits_16_and_inst14_in1 = {magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out};
	coreir_and #(.width(16)) magma_Bits_16_and_inst14(
		.in0(a),
		.in1(magma_Bits_16_and_inst14_in1),
		.out(magma_Bits_16_and_inst14_out)
	);
	wire [15:0] magma_Bits_16_and_inst15_in1;
	assign magma_Bits_16_and_inst15_in1 = {magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out, magma_Bits_8_eq_inst30_out};
	coreir_and #(.width(16)) magma_Bits_16_and_inst15(
		.in0(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(magma_Bits_16_and_inst15_in1),
		.out(magma_Bits_16_and_inst15_out)
	);
	wire [15:0] magma_Bits_16_and_inst16_in1;
	assign magma_Bits_16_and_inst16_in1 = {magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out};
	coreir_and #(.width(16)) magma_Bits_16_and_inst16(
		.in0(a),
		.in1(magma_Bits_16_and_inst16_in1),
		.out(magma_Bits_16_and_inst16_out)
	);
	wire [15:0] magma_Bits_16_and_inst17_in1;
	assign magma_Bits_16_and_inst17_in1 = {magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out, magma_Bit_or_inst7_out};
	coreir_and #(.width(16)) magma_Bits_16_and_inst17(
		.in0(Mux2xBits16_inst12$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(magma_Bits_16_and_inst17_in1),
		.out(magma_Bits_16_and_inst17_out)
	);
	coreir_and #(.width(16)) magma_Bits_16_and_inst2(
		.in0(a),
		.in1(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.out(magma_Bits_16_and_inst2_out)
	);
	coreir_and #(.width(16)) magma_Bits_16_and_inst3(
		.in0(a),
		.in1(const_127_16_out),
		.out(magma_Bits_16_and_inst3_out)
	);
	coreir_and #(.width(16)) magma_Bits_16_and_inst4(
		.in0(a),
		.in1(const_32768_16_out),
		.out(magma_Bits_16_and_inst4_out)
	);
	coreir_and #(.width(16)) magma_Bits_16_and_inst5(
		.in0(a),
		.in1(const_127_16_out),
		.out(magma_Bits_16_and_inst5_out)
	);
	coreir_and #(.width(16)) magma_Bits_16_and_inst6(
		.in0(a),
		.in1(const_32768_16_out),
		.out(magma_Bits_16_and_inst6_out)
	);
	coreir_and #(.width(16)) magma_Bits_16_and_inst7(
		.in0(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_32768_16_out),
		.out(magma_Bits_16_and_inst7_out)
	);
	coreir_and #(.width(16)) magma_Bits_16_and_inst8(
		.in0(a),
		.in1(const_127_16_out),
		.out(magma_Bits_16_and_inst8_out)
	);
	coreir_and #(.width(16)) magma_Bits_16_and_inst9(
		.in0(a),
		.in1(const_32768_16_out),
		.out(magma_Bits_16_and_inst9_out)
	);
	coreir_eq #(.width(16)) magma_Bits_16_eq_inst0(
		.in0(magma_Bits_16_and_inst9_out),
		.in1(const_32768_16_out),
		.out(magma_Bits_16_eq_inst0_out)
	);
	coreir_eq #(.width(16)) magma_Bits_16_eq_inst1(
		.in0(magma_Bits_16_and_inst11_out),
		.in1(const_32768_16_out),
		.out(magma_Bits_16_eq_inst1_out)
	);
	coreir_lshr #(.width(16)) magma_Bits_16_lshr_inst0(
		.in0(Mux2xBits16_inst5$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_8_16_out),
		.out(magma_Bits_16_lshr_inst0_out)
	);
	wire [15:0] magma_Bits_16_lshr_inst1_in1;
	assign magma_Bits_16_lshr_inst1_in1 = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, magma_SInt_9_neg_inst1_out[8:0]};
	coreir_lshr #(.width(16)) magma_Bits_16_lshr_inst1(
		.in0(magma_Bits_16_or_inst9_out),
		.in1(magma_Bits_16_lshr_inst1_in1),
		.out(magma_Bits_16_lshr_inst1_out)
	);
	coreir_not #(.width(16)) magma_Bits_16_not_inst0(
		.in(b),
		.out(magma_Bits_16_not_inst0_out)
	);
	coreir_or #(.width(16)) magma_Bits_16_or_inst0(
		.in0(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(magma_Bits_16_and_inst1_out),
		.out(magma_Bits_16_or_inst0_out)
	);
	coreir_or #(.width(16)) magma_Bits_16_or_inst1(
		.in0(magma_Bits_16_or_inst0_out),
		.in1(Mux2xBits16_inst6$coreir_commonlib_mux2x16_inst0$_join_out),
		.out(magma_Bits_16_or_inst1_out)
	);
	coreir_or #(.width(16)) magma_Bits_16_or_inst2(
		.in0(a),
		.in1(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.out(magma_Bits_16_or_inst2_out)
	);
	coreir_or #(.width(16)) magma_Bits_16_or_inst3(
		.in0(magma_Bits_16_and_inst4_out),
		.in1(magma_Bits_16_shl_inst3_out),
		.out(magma_Bits_16_or_inst3_out)
	);
	coreir_or #(.width(16)) magma_Bits_16_or_inst4(
		.in0(magma_Bits_16_or_inst3_out),
		.in1(magma_Bits_16_and_inst5_out),
		.out(magma_Bits_16_or_inst4_out)
	);
	coreir_or #(.width(16)) magma_Bits_16_or_inst5(
		.in0(magma_Bits_16_and_inst6_out),
		.in1(magma_Bits_16_and_inst7_out),
		.out(magma_Bits_16_or_inst5_out)
	);
	coreir_or #(.width(16)) magma_Bits_16_or_inst6(
		.in0(magma_Bits_16_or_inst5_out),
		.in1(magma_Bits_16_shl_inst4_out),
		.out(magma_Bits_16_or_inst6_out)
	);
	coreir_or #(.width(16)) magma_Bits_16_or_inst7(
		.in0(magma_Bits_16_or_inst6_out),
		.in1(magma_Bits_16_and_inst8_out),
		.out(magma_Bits_16_or_inst7_out)
	);
	coreir_or #(.width(16)) magma_Bits_16_or_inst8(
		.in0(magma_Bits_16_and_inst10_out),
		.in1(const_128_16_out),
		.out(magma_Bits_16_or_inst8_out)
	);
	coreir_or #(.width(16)) magma_Bits_16_or_inst9(
		.in0(magma_Bits_16_and_inst12_out),
		.in1(const_128_16_out),
		.out(magma_Bits_16_or_inst9_out)
	);
	coreir_shl #(.width(16)) magma_Bits_16_shl_inst0(
		.in0(magma_SInt_16_add_inst0_out),
		.in1(const_7_16_out),
		.out(magma_Bits_16_shl_inst0_out)
	);
	coreir_shl #(.width(16)) magma_Bits_16_shl_inst1(
		.in0(a),
		.in1(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.out(magma_Bits_16_shl_inst1_out)
	);
	coreir_shl #(.width(16)) magma_Bits_16_shl_inst2(
		.in0(const_1_16_out),
		.in1(const_15_16_out),
		.out(magma_Bits_16_shl_inst2_out)
	);
	wire [15:0] magma_Bits_16_shl_inst3_in0;
	assign magma_Bits_16_shl_inst3_in0 = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, magma_UInt_8_add_inst0_out[7:0]};
	coreir_shl #(.width(16)) magma_Bits_16_shl_inst3(
		.in0(magma_Bits_16_shl_inst3_in0),
		.in1(const_7_16_out),
		.out(magma_Bits_16_shl_inst3_out)
	);
	wire [15:0] magma_Bits_16_shl_inst4_in0;
	assign magma_Bits_16_shl_inst4_in0 = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, magma_UInt_8_add_inst1_out[7:0]};
	coreir_shl #(.width(16)) magma_Bits_16_shl_inst4(
		.in0(magma_Bits_16_shl_inst4_in0),
		.in1(const_7_16_out),
		.out(magma_Bits_16_shl_inst4_out)
	);
	wire [15:0] magma_Bits_16_shl_inst5_in1;
	assign magma_Bits_16_shl_inst5_in1 = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, magma_SInt_9_sub_inst2_out[8:0]};
	coreir_shl #(.width(16)) magma_Bits_16_shl_inst5(
		.in0(magma_Bits_16_or_inst9_out),
		.in1(magma_Bits_16_shl_inst5_in1),
		.out(magma_Bits_16_shl_inst5_out)
	);
	coreir_xor #(.width(16)) magma_Bits_16_xor_inst0(
		.in0(a),
		.in1(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.out(magma_Bits_16_xor_inst0_out)
	);
	coreir_xor #(.width(16)) magma_Bits_16_xor_inst1(
		.in0(magma_Bits_16_shl_inst2_out),
		.in1(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.out(magma_Bits_16_xor_inst1_out)
	);
	coreir_eq #(.width(1)) magma_Bits_1_eq_inst0(
		.in0(signed_),
		.in1(const_1_1_out),
		.out(magma_Bits_1_eq_inst0_out)
	);
	coreir_eq #(.width(1)) magma_Bits_1_eq_inst1(
		.in0(signed_),
		.in1(const_1_1_out),
		.out(magma_Bits_1_eq_inst1_out)
	);
	coreir_lshr #(.width(23)) magma_Bits_23_lshr_inst0(
		.in0(Mux2xBits23_inst0$coreir_commonlib_mux2x23_inst0$_join_out),
		.in1(const_7_23_out),
		.out(magma_Bits_23_lshr_inst0_out)
	);
	wire [22:0] magma_Bits_23_shl_inst0_in0;
	assign magma_Bits_23_shl_inst0_in0 = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, magma_Bits_16_or_inst8_out[15:0]};
	wire [22:0] magma_Bits_23_shl_inst0_in1;
	assign magma_Bits_23_shl_inst0_in1 = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, magma_SInt_9_sub_inst1_out[8:0]};
	coreir_shl #(.width(23)) magma_Bits_23_shl_inst0(
		.in0(magma_Bits_23_shl_inst0_in0),
		.in1(magma_Bits_23_shl_inst0_in1),
		.out(magma_Bits_23_shl_inst0_out)
	);
	coreir_eq #(.width(7)) magma_Bits_7_eq_inst0(
		.in0(a[6:0]),
		.in1(const_0_7_out),
		.out(magma_Bits_7_eq_inst0_out)
	);
	coreir_eq #(.width(7)) magma_Bits_7_eq_inst1(
		.in0(b[6:0]),
		.in1(const_0_7_out),
		.out(magma_Bits_7_eq_inst1_out)
	);
	coreir_eq #(.width(7)) magma_Bits_7_eq_inst2(
		.in0(Mux2xBits16_inst70_O_out[6:0]),
		.in1(const_0_7_out),
		.out(magma_Bits_7_eq_inst2_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst0(
		.in0(a[14:7]),
		.in1(const_255_8_out),
		.out(magma_Bits_8_eq_inst0_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst1(
		.in0(b[14:7]),
		.in1(const_255_8_out),
		.out(magma_Bits_8_eq_inst1_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst10(
		.in0(alu),
		.in1(const_1_8_out),
		.out(magma_Bits_8_eq_inst10_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst11(
		.in0(alu),
		.in1(const_2_8_out),
		.out(magma_Bits_8_eq_inst11_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst12(
		.in0(alu),
		.in1(const_6_8_out),
		.out(magma_Bits_8_eq_inst12_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst13(
		.in0(alu),
		.in1(const_11_8_out),
		.out(magma_Bits_8_eq_inst13_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst14(
		.in0(alu),
		.in1(const_12_8_out),
		.out(magma_Bits_8_eq_inst14_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst15(
		.in0(alu),
		.in1(const_13_8_out),
		.out(magma_Bits_8_eq_inst15_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst16(
		.in0(alu),
		.in1(const_4_8_out),
		.out(magma_Bits_8_eq_inst16_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst17(
		.in0(alu),
		.in1(const_5_8_out),
		.out(magma_Bits_8_eq_inst17_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst18(
		.in0(alu),
		.in1(const_3_8_out),
		.out(magma_Bits_8_eq_inst18_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst19(
		.in0(alu),
		.in1(const_8_8_out),
		.out(magma_Bits_8_eq_inst19_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst2(
		.in0(alu),
		.in1(const_149_8_out),
		.out(magma_Bits_8_eq_inst2_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst20(
		.in0(alu),
		.in1(const_19_8_out),
		.out(magma_Bits_8_eq_inst20_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst21(
		.in0(alu),
		.in1(const_18_8_out),
		.out(magma_Bits_8_eq_inst21_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst22(
		.in0(alu),
		.in1(const_20_8_out),
		.out(magma_Bits_8_eq_inst22_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst23(
		.in0(alu),
		.in1(const_15_8_out),
		.out(magma_Bits_8_eq_inst23_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst24(
		.in0(alu),
		.in1(const_17_8_out),
		.out(magma_Bits_8_eq_inst24_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst25(
		.in0(alu),
		.in1(const_22_8_out),
		.out(magma_Bits_8_eq_inst25_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst26(
		.in0(alu),
		.in1(const_23_8_out),
		.out(magma_Bits_8_eq_inst26_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst27(
		.in0(alu),
		.in1(const_24_8_out),
		.out(magma_Bits_8_eq_inst27_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst28(
		.in0(alu),
		.in1(const_23_8_out),
		.out(magma_Bits_8_eq_inst28_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst29(
		.in0(alu),
		.in1(const_24_8_out),
		.out(magma_Bits_8_eq_inst29_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst3(
		.in0(alu),
		.in1(const_152_8_out),
		.out(magma_Bits_8_eq_inst3_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst30(
		.in0(alu),
		.in1(const_25_8_out),
		.out(magma_Bits_8_eq_inst30_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst31(
		.in0(alu),
		.in1(const_146_8_out),
		.out(magma_Bits_8_eq_inst31_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst32(
		.in0(alu),
		.in1(const_147_8_out),
		.out(magma_Bits_8_eq_inst32_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst33(
		.in0(alu),
		.in1(const_148_8_out),
		.out(magma_Bits_8_eq_inst33_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst34(
		.in0(alu),
		.in1(const_149_8_out),
		.out(magma_Bits_8_eq_inst34_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst35(
		.in0(alu),
		.in1(const_150_8_out),
		.out(magma_Bits_8_eq_inst35_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst36(
		.in0(alu),
		.in1(const_151_8_out),
		.out(magma_Bits_8_eq_inst36_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst37(
		.in0(alu),
		.in1(const_23_8_out),
		.out(magma_Bits_8_eq_inst37_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst38(
		.in0(alu),
		.in1(const_22_8_out),
		.out(magma_Bits_8_eq_inst38_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst39(
		.in0(alu),
		.in1(const_25_8_out),
		.out(magma_Bits_8_eq_inst39_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst4(
		.in0(alu),
		.in1(const_1_8_out),
		.out(magma_Bits_8_eq_inst4_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst40(
		.in0(alu),
		.in1(const_24_8_out),
		.out(magma_Bits_8_eq_inst40_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst41(
		.in0(Mux2xBits16_inst70_O_out[14:7]),
		.in1(const_0_8_out),
		.out(magma_Bits_8_eq_inst41_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst42(
		.in0(alu),
		.in1(const_24_8_out),
		.out(magma_Bits_8_eq_inst42_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst5(
		.in0(alu),
		.in1(const_6_8_out),
		.out(magma_Bits_8_eq_inst5_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst6(
		.in0(alu),
		.in1(const_1_8_out),
		.out(magma_Bits_8_eq_inst6_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst7(
		.in0(alu),
		.in1(const_2_8_out),
		.out(magma_Bits_8_eq_inst7_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst8(
		.in0(alu),
		.in1(const_6_8_out),
		.out(magma_Bits_8_eq_inst8_out)
	);
	coreir_eq #(.width(8)) magma_Bits_8_eq_inst9(
		.in0(alu),
		.in1(const_0_8_out),
		.out(magma_Bits_8_eq_inst9_out)
	);
	coreir_add #(.width(16)) magma_SInt_16_add_inst0(
		.in0(Mux2xSInt16_inst27$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_127_16_out),
		.out(magma_SInt_16_add_inst0_out)
	);
	coreir_and #(.width(16)) magma_SInt_16_and_inst0(
		.in0(magma_SInt_16_shl_inst0_out),
		.in1(Mux2xSInt16_inst24$coreir_commonlib_mux2x16_inst0$_join_out),
		.out(magma_SInt_16_and_inst0_out)
	);
	coreir_ashr #(.width(16)) magma_SInt_16_ashr_inst0(
		.in0(a),
		.in1(b),
		.out(magma_SInt_16_ashr_inst0_out)
	);
	coreir_eq #(.width(16)) magma_SInt_16_eq_inst0(
		.in0(const_0_16_out),
		.in1(Mux2xBits16_inst70$coreir_commonlib_mux2x16_inst0$_join_out),
		.out(magma_SInt_16_eq_inst0_out)
	);
	coreir_neg #(.width(16)) magma_SInt_16_neg_inst0(
		.in(a),
		.out(magma_SInt_16_neg_inst0_out)
	);
	coreir_neg #(.width(16)) magma_SInt_16_neg_inst1(
		.in(a),
		.out(magma_SInt_16_neg_inst1_out)
	);
	coreir_neg #(.width(16)) magma_SInt_16_neg_inst2(
		.in(magma_Bits_23_lshr_inst0_out[15:0]),
		.out(magma_SInt_16_neg_inst2_out)
	);
	coreir_neg #(.width(16)) magma_SInt_16_neg_inst3(
		.in(magma_Bits_16_and_inst13_out),
		.out(magma_SInt_16_neg_inst3_out)
	);
	coreir_sge #(.width(16)) magma_SInt_16_sge_inst0(
		.in0(a),
		.in1(b),
		.out(magma_SInt_16_sge_inst0_out)
	);
	coreir_sge #(.width(16)) magma_SInt_16_sge_inst1(
		.in0(a),
		.in1(const_0_16_out),
		.out(magma_SInt_16_sge_inst1_out)
	);
	coreir_sge #(.width(16)) magma_SInt_16_sge_inst2(
		.in0(Mux2xSInt16_inst27$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(const_0_16_out),
		.out(magma_SInt_16_sge_inst2_out)
	);
	coreir_shl #(.width(16)) magma_SInt_16_shl_inst0(
		.in0(Mux2xSInt16_inst25$coreir_commonlib_mux2x16_inst0$_join_out),
		.in1(Mux2xSInt16_inst26$coreir_commonlib_mux2x16_inst0$_join_out),
		.out(magma_SInt_16_shl_inst0_out)
	);
	coreir_sle #(.width(16)) magma_SInt_16_sle_inst0(
		.in0(a),
		.in1(b),
		.out(magma_SInt_16_sle_inst0_out)
	);
	coreir_sub #(.width(16)) magma_SInt_16_sub_inst0(
		.in0(const_7_16_out),
		.in1(Mux2xSInt16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
		.out(magma_SInt_16_sub_inst0_out)
	);
	coreir_sub #(.width(16)) magma_SInt_16_sub_inst1(
		.in0(const_15_16_out),
		.in1(Mux2xSInt16_inst23$coreir_commonlib_mux2x16_inst0$_join_out),
		.out(magma_SInt_16_sub_inst1_out)
	);
	coreir_neg #(.width(9)) magma_SInt_9_neg_inst0(
		.in(magma_SInt_9_sub_inst0_out),
		.out(magma_SInt_9_neg_inst0_out)
	);
	coreir_neg #(.width(9)) magma_SInt_9_neg_inst1(
		.in(magma_SInt_9_sub_inst2_out),
		.out(magma_SInt_9_neg_inst1_out)
	);
	coreir_slt #(.width(9)) magma_SInt_9_slt_inst0(
		.in0(magma_SInt_9_sub_inst0_out),
		.in1(const_0_9_out),
		.out(magma_SInt_9_slt_inst0_out)
	);
	coreir_slt #(.width(9)) magma_SInt_9_slt_inst1(
		.in0(magma_SInt_9_sub_inst1_out),
		.in1(const_0_9_out),
		.out(magma_SInt_9_slt_inst1_out)
	);
	coreir_slt #(.width(9)) magma_SInt_9_slt_inst2(
		.in0(magma_SInt_9_sub_inst2_out),
		.in1(const_0_9_out),
		.out(magma_SInt_9_slt_inst2_out)
	);
	wire [8:0] magma_SInt_9_sub_inst0_in0;
	assign magma_SInt_9_sub_inst0_in0 = {bit_const_0_None_out, a[14:7]};
	coreir_sub #(.width(9)) magma_SInt_9_sub_inst0(
		.in0(magma_SInt_9_sub_inst0_in0),
		.in1(const_127_9_out),
		.out(magma_SInt_9_sub_inst0_out)
	);
	wire [8:0] magma_SInt_9_sub_inst1_in0;
	assign magma_SInt_9_sub_inst1_in0 = {bit_const_0_None_out, a[14:7]};
	coreir_sub #(.width(9)) magma_SInt_9_sub_inst1(
		.in0(magma_SInt_9_sub_inst1_in0),
		.in1(const_127_9_out),
		.out(magma_SInt_9_sub_inst1_out)
	);
	wire [8:0] magma_SInt_9_sub_inst2_in0;
	assign magma_SInt_9_sub_inst2_in0 = {bit_const_0_None_out, a[14:7]};
	coreir_sub #(.width(9)) magma_SInt_9_sub_inst2(
		.in0(magma_SInt_9_sub_inst2_in0),
		.in1(const_127_9_out),
		.out(magma_SInt_9_sub_inst2_out)
	);
	coreir_lshr #(.width(16)) magma_UInt_16_lshr_inst0(
		.in0(a),
		.in1(b),
		.out(magma_UInt_16_lshr_inst0_out)
	);
	coreir_uge #(.width(16)) magma_UInt_16_uge_inst0(
		.in0(a),
		.in1(b),
		.out(magma_UInt_16_uge_inst0_out)
	);
	coreir_ule #(.width(16)) magma_UInt_16_ule_inst0(
		.in0(a),
		.in1(b),
		.out(magma_UInt_16_ule_inst0_out)
	);
	wire [16:0] magma_UInt_17_add_inst0_in0;
	assign magma_UInt_17_add_inst0_in0 = {bit_const_0_None_out, a[15:0]};
	wire [16:0] magma_UInt_17_add_inst0_in1;
	assign magma_UInt_17_add_inst0_in1 = {bit_const_0_None_out, Mux2xBits16_inst7_O_out[15:0]};
	coreir_add #(.width(17)) magma_UInt_17_add_inst0(
		.in0(magma_UInt_17_add_inst0_in0),
		.in1(magma_UInt_17_add_inst0_in1),
		.out(magma_UInt_17_add_inst0_out)
	);
	wire [16:0] magma_UInt_17_add_inst1_in1;
	assign magma_UInt_17_add_inst1_in1 = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out[0]};
	coreir_add #(.width(17)) magma_UInt_17_add_inst1(
		.in0(magma_UInt_17_add_inst0_out),
		.in1(magma_UInt_17_add_inst1_in1),
		.out(magma_UInt_17_add_inst1_out)
	);
	wire [31:0] magma_UInt_32_and_inst0_in1;
	assign magma_UInt_32_and_inst0_in1 = {magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out};
	coreir_and #(.width(32)) magma_UInt_32_and_inst0(
		.in0(Mux2xUInt32_inst0$coreir_commonlib_mux2x32_inst0$_join_out),
		.in1(magma_UInt_32_and_inst0_in1),
		.out(magma_UInt_32_and_inst0_out)
	);
	wire [31:0] magma_UInt_32_and_inst1_in1;
	assign magma_UInt_32_and_inst1_in1 = {magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out, magma_Bit_or_inst13_out};
	coreir_and #(.width(32)) magma_UInt_32_and_inst1(
		.in0(Mux2xUInt32_inst1$coreir_commonlib_mux2x32_inst0$_join_out),
		.in1(magma_UInt_32_and_inst1_in1),
		.out(magma_UInt_32_and_inst1_out)
	);
	coreir_mul #(.width(32)) magma_UInt_32_mul_inst0(
		.in0(magma_UInt_32_and_inst0_out),
		.in1(magma_UInt_32_and_inst1_out),
		.out(magma_UInt_32_mul_inst0_out)
	);
	coreir_add #(.width(8)) magma_UInt_8_add_inst0(
		.in0(a[14:7]),
		.in1(Mux2xBits16_inst7_O_out[7:0]),
		.out(magma_UInt_8_add_inst0_out)
	);
	coreir_add #(.width(8)) magma_UInt_8_add_inst1(
		.in0(magma_UInt_8_sub_inst0_out),
		.in1(const_127_8_out),
		.out(magma_UInt_8_add_inst1_out)
	);
	coreir_sub #(.width(8)) magma_UInt_8_sub_inst0(
		.in0(a[14:7]),
		.in1(Mux2xBits16_inst7_O_out[14:7]),
		.out(magma_UInt_8_sub_inst0_out)
	);
	coreir_ugt #(.width(8)) magma_UInt_8_ugt_inst0(
		.in0(a[14:7]),
		.in1(const_142_8_out),
		.out(magma_UInt_8_ugt_inst0_out)
	);
	wire [8:0] magma_UInt_9_add_inst0_in0;
	assign magma_UInt_9_add_inst0_in0 = {bit_const_0_None_out, a[14:7]};
	coreir_add #(.width(9)) magma_UInt_9_add_inst0(
		.in0(magma_UInt_9_add_inst0_in0),
		.in1(Mux2xBits16_inst7_O_out[8:0]),
		.out(magma_UInt_9_add_inst0_out)
	);
	coreir_ugt #(.width(9)) magma_UInt_9_ugt_inst0(
		.in0(magma_UInt_9_add_inst0_out),
		.in1(const_255_9_out),
		.out(magma_UInt_9_ugt_inst0_out)
	);
	assign O0 = Mux2xBits16_inst70$coreir_commonlib_mux2x16_inst0$_join_out;
	assign O1 = Mux2xBit_inst49$coreir_commonlib_mux2x1_inst0$_join_out[0];
	assign O2 = Mux2xBit_inst52$coreir_commonlib_mux2x1_inst0$_join_out[0];
	assign O3 = Mux2xBits16_inst70_O_out[15];
	assign O4 = Mux2xBit_inst47$coreir_commonlib_mux2x1_inst0$_join_out[0];
	assign O5 = Mux2xBit_inst48$coreir_commonlib_mux2x1_inst0$_join_out[0];
endmodule
module PE (
	inst,
	data0,
	data1,
	bit0,
	bit1,
	bit2,
	clk_en,
	config_addr,
	config_data,
	config_en,
	O0,
	O1,
	O2,
	CLK,
	ASYNCRESET
);
	input [66:0] inst;
	input [15:0] data0;
	input [15:0] data1;
	input bit0;
	input bit1;
	input bit2;
	input clk_en;
	input [7:0] config_addr;
	input [31:0] config_data;
	input config_en;
	output [15:0] O0;
	output O1;
	output [31:0] O2;
	input CLK;
	input ASYNCRESET;
	wire [15:0] ALU_inst0_O0;
	wire ALU_inst0_O1;
	wire ALU_inst0_O2;
	wire ALU_inst0_O3;
	wire ALU_inst0_O4;
	wire ALU_inst0_O5;
	wire Cond_inst0_O;
	wire LUT_inst0_O;
	wire [0:0] Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBits1_inst1$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [0:0] Mux2xBits1_inst2$coreir_commonlib_mux2x1_inst0$_join_out;
	wire [31:0] Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
	wire [31:0] Mux2xBits32_inst0_I0_in;
	wire [15:0] RegisterMode_inst0_O0;
	wire [15:0] RegisterMode_inst0_O1;
	wire [15:0] RegisterMode_inst1_O0;
	wire [15:0] RegisterMode_inst1_O1;
	wire RegisterMode_inst2_O0;
	wire RegisterMode_inst2_O1;
	wire RegisterMode_inst3_O0;
	wire RegisterMode_inst3_O1;
	wire RegisterMode_inst4_O0;
	wire RegisterMode_inst4_O1;
	wire bit_const_0_None_out;
	wire [0:0] const_0_1_out;
	wire [0:0] const_1_1_out;
	wire [2:0] const_3_3_out;
	wire [2:0] const_4_3_out;
	wire magma_Bit_and_inst0_out;
	wire magma_Bit_and_inst1_out;
	wire magma_Bits_3_eq_inst0_out;
	wire magma_Bits_3_eq_inst1_out;
	ALU ALU_inst0(
		.alu(inst[7:0]),
		.signed_(inst[8]),
		.a(RegisterMode_inst0_O0),
		.b(RegisterMode_inst1_O0),
		.d(RegisterMode_inst2_O0),
		.O0(ALU_inst0_O0),
		.O1(ALU_inst0_O1),
		.O2(ALU_inst0_O2),
		.O3(ALU_inst0_O3),
		.O4(ALU_inst0_O4),
		.O5(ALU_inst0_O5),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	Cond Cond_inst0(
		.code(inst[21:17]),
		.alu(ALU_inst0_O1),
		.lut(LUT_inst0_O),
		.Z(ALU_inst0_O2),
		.N(ALU_inst0_O3),
		.C(ALU_inst0_O4),
		.V(ALU_inst0_O5),
		.O(Cond_inst0_O),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	LUT LUT_inst0(
		.lut(inst[16:9]),
		.bit0(RegisterMode_inst2_O0),
		.bit1(RegisterMode_inst3_O0),
		.bit2(RegisterMode_inst4_O0),
		.O(LUT_inst0_O),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	coreir_mux #(.width(1)) Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
		.in0(const_0_1_out),
		.in1(const_1_1_out),
		.sel(RegisterMode_inst2_O1),
		.out(Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBits1_inst1$coreir_commonlib_mux2x1_inst0$_join(
		.in0(const_0_1_out),
		.in1(const_1_1_out),
		.sel(RegisterMode_inst3_O1),
		.out(Mux2xBits1_inst1$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	coreir_mux #(.width(1)) Mux2xBits1_inst2$coreir_commonlib_mux2x1_inst0$_join(
		.in0(const_0_1_out),
		.in1(const_1_1_out),
		.sel(RegisterMode_inst4_O1),
		.out(Mux2xBits1_inst2$coreir_commonlib_mux2x1_inst0$_join_out)
	);
	wire [31:0] Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_in1;
	assign Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_in1 = {bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, bit_const_0_None_out, Mux2xBits1_inst2$coreir_commonlib_mux2x1_inst0$_join_out[0], Mux2xBits1_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0], Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]};
	coreir_mux #(.width(32)) Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join(
		.in0(Mux2xBits32_inst0_I0_in),
		.in1(Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_in1),
		.sel(magma_Bits_3_eq_inst1_out),
		.out(Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out)
	);
	wire [31:0] Mux2xBits32_inst0_I0_out;
	assign Mux2xBits32_inst0_I0_out = {RegisterMode_inst1_O1[15:0], RegisterMode_inst0_O1[15:0]};
	mantle_wire__typeBitIn32 Mux2xBits32_inst0_I0(
		.in(Mux2xBits32_inst0_I0_in),
		.out(Mux2xBits32_inst0_I0_out)
	);
	RegisterMode RegisterMode_inst0(
		.mode(inst[23:22]),
		.const_(inst[39:24]),
		.value(data0),
		.clk_en(clk_en),
		.config_we(magma_Bit_and_inst0_out),
		.config_data(config_data[15:0]),
		.O0(RegisterMode_inst0_O0),
		.O1(RegisterMode_inst0_O1),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	RegisterMode RegisterMode_inst1(
		.mode(inst[41:40]),
		.const_(inst[57:42]),
		.value(data1),
		.clk_en(clk_en),
		.config_we(magma_Bit_and_inst0_out),
		.config_data(config_data[31:16]),
		.O0(RegisterMode_inst1_O0),
		.O1(RegisterMode_inst1_O1),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	RegisterMode_unq1 RegisterMode_inst2(
		.mode(inst[59:58]),
		.const_(inst[60]),
		.value(bit0),
		.clk_en(clk_en),
		.config_we(magma_Bit_and_inst1_out),
		.config_data(config_data[0]),
		.O0(RegisterMode_inst2_O0),
		.O1(RegisterMode_inst2_O1),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	RegisterMode_unq1 RegisterMode_inst3(
		.mode(inst[62:61]),
		.const_(inst[63]),
		.value(bit1),
		.clk_en(clk_en),
		.config_we(magma_Bit_and_inst1_out),
		.config_data(config_data[1]),
		.O0(RegisterMode_inst3_O0),
		.O1(RegisterMode_inst3_O1),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	RegisterMode_unq1 RegisterMode_inst4(
		.mode(inst[65:64]),
		.const_(inst[66]),
		.value(bit2),
		.clk_en(clk_en),
		.config_we(magma_Bit_and_inst1_out),
		.config_data(config_data[2]),
		.O0(RegisterMode_inst4_O0),
		.O1(RegisterMode_inst4_O1),
		.CLK(CLK),
		.ASYNCRESET(ASYNCRESET)
	);
	corebit_const #(.value(1'b0)) bit_const_0_None(.out(bit_const_0_None_out));
	coreir_const #(
		.value(1'h0),
		.width(1)
	) const_0_1(.out(const_0_1_out));
	coreir_const #(
		.value(1'h1),
		.width(1)
	) const_1_1(.out(const_1_1_out));
	coreir_const #(
		.value(3'h3),
		.width(3)
	) const_3_3(.out(const_3_3_out));
	coreir_const #(
		.value(3'h4),
		.width(3)
	) const_4_3(.out(const_4_3_out));
	corebit_and magma_Bit_and_inst0(
		.in0(magma_Bits_3_eq_inst0_out),
		.in1(config_en),
		.out(magma_Bit_and_inst0_out)
	);
	corebit_and magma_Bit_and_inst1(
		.in0(magma_Bits_3_eq_inst1_out),
		.in1(config_en),
		.out(magma_Bit_and_inst1_out)
	);
	coreir_eq #(.width(3)) magma_Bits_3_eq_inst0(
		.in0(config_addr[2:0]),
		.in1(const_3_3_out),
		.out(magma_Bits_3_eq_inst0_out)
	);
	coreir_eq #(.width(3)) magma_Bits_3_eq_inst1(
		.in0(config_addr[2:0]),
		.in1(const_4_3_out),
		.out(magma_Bits_3_eq_inst1_out)
	);
	assign O0 = ALU_inst0_O0;
	assign O1 = Cond_inst0_O;
	assign O2 = Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
endmodule
module PE_unq1 (
	alu_res,
	bit0,
	bit1,
	bit2,
	clk,
	config_config_addr,
	config_config_data,
	config_read,
	config_write,
	data0,
	data1,
	read_config_data,
	res_p,
	reset,
	stall
);
	output [15:0] alu_res;
	input [0:0] bit0;
	input [0:0] bit1;
	input [0:0] bit2;
	input clk;
	input [7:0] config_config_addr;
	input [31:0] config_config_data;
	input [0:0] config_read;
	input [0:0] config_write;
	input [15:0] data0;
	input [15:0] data1;
	output [31:0] read_config_data;
	output [0:0] res_p;
	input reset;
	input [0:0] stall;
	wire [0:0] Invert1_inst0_out;
	wire [31:0] MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0_out;
	wire [1:0] MuxWrapper_3_32_inst0_S_in;
	wire [15:0] WrappedPE_inst0$PE_inst0_O0;
	wire WrappedPE_inst0$PE_inst0_O1;
	wire [31:0] WrappedPE_inst0$PE_inst0_O2;
	wire [66:0] WrappedPE_inst0_inst_in;
	wire bit_const_0_None_out;
	wire [31:0] config_reg_0_O;
	wire [31:0] config_reg_1_O;
	wire [31:0] config_reg_2_O;
	wire [31:0] inst_0_inst0_O;
	wire [31:0] inst_1_inst0_O;
	wire [31:0] inst_2_inst0_O;
	wire [7:0] self_config_config_addr_out;
	coreir_not #(.width(1)) Invert1_inst0(
		.in(stall),
		.out(Invert1_inst0_out)
	);
	commonlib_muxn__N3__width32 MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0(
		.in_data_0(config_reg_0_O),
		.in_data_1(config_reg_1_O),
		.in_data_2(config_reg_2_O),
		.in_sel(MuxWrapper_3_32_inst0_S_in),
		.out(MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0_out)
	);
	mantle_wire__typeBitIn2 MuxWrapper_3_32_inst0_S(
		.in(MuxWrapper_3_32_inst0_S_in),
		.out(self_config_config_addr_out[1:0])
	);
	PE WrappedPE_inst0$PE_inst0(
		.inst(WrappedPE_inst0_inst_in),
		.data0(data0),
		.data1(data1),
		.bit0(bit0[0]),
		.bit1(bit1[0]),
		.bit2(bit2[0]),
		.clk_en(Invert1_inst0_out[0]),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(bit_const_0_None_out),
		.O0(WrappedPE_inst0$PE_inst0_O0),
		.O1(WrappedPE_inst0$PE_inst0_O1),
		.O2(WrappedPE_inst0$PE_inst0_O2),
		.CLK(clk),
		.ASYNCRESET(reset)
	);
	wire [66:0] WrappedPE_inst0_inst_out;
	assign WrappedPE_inst0_inst_out = {inst_2_inst0_O[2:0], inst_1_inst0_O[31:0], inst_0_inst0_O[31:0]};
	mantle_wire__typeBitIn67 WrappedPE_inst0_inst(
		.in(WrappedPE_inst0_inst_in),
		.out(WrappedPE_inst0_inst_out)
	);
	corebit_const #(.value(1'b0)) bit_const_0_None(.out(bit_const_0_None_out));
	ConfigRegister_32_8_32_0 config_reg_0(
		.clk(clk),
		.reset(reset),
		.O(config_reg_0_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_1 config_reg_1(
		.clk(clk),
		.reset(reset),
		.O(config_reg_1_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	ConfigRegister_32_8_32_2 config_reg_2(
		.clk(clk),
		.reset(reset),
		.O(config_reg_2_O),
		.config_addr(config_config_addr),
		.config_data(config_config_data),
		.config_en(config_write[0])
	);
	inst_0 inst_0_inst0(
		.I(config_reg_0_O),
		.O(inst_0_inst0_O)
	);
	inst_1 inst_1_inst0(
		.I(config_reg_1_O),
		.O(inst_1_inst0_O)
	);
	inst_2 inst_2_inst0(
		.I(config_reg_2_O),
		.O(inst_2_inst0_O)
	);
	mantle_wire__typeBit8 self_config_config_addr(
		.in(config_config_addr),
		.out(self_config_config_addr_out)
	);
	assign alu_res = WrappedPE_inst0$PE_inst0_O0;
	assign read_config_data = MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0_out;
	assign res_p = WrappedPE_inst0$PE_inst0_O1;
endmodule
module Tile_PE (
	SB_T0_EAST_SB_IN_B1,
	SB_T0_EAST_SB_IN_B16,
	SB_T0_EAST_SB_OUT_B1,
	SB_T0_EAST_SB_OUT_B16,
	SB_T0_NORTH_SB_IN_B1,
	SB_T0_NORTH_SB_IN_B16,
	SB_T0_NORTH_SB_OUT_B1,
	SB_T0_NORTH_SB_OUT_B16,
	SB_T0_SOUTH_SB_IN_B1,
	SB_T0_SOUTH_SB_IN_B16,
	SB_T0_SOUTH_SB_OUT_B1,
	SB_T0_SOUTH_SB_OUT_B16,
	SB_T0_WEST_SB_IN_B1,
	SB_T0_WEST_SB_IN_B16,
	SB_T0_WEST_SB_OUT_B1,
	SB_T0_WEST_SB_OUT_B16,
	SB_T1_EAST_SB_IN_B1,
	SB_T1_EAST_SB_IN_B16,
	SB_T1_EAST_SB_OUT_B1,
	SB_T1_EAST_SB_OUT_B16,
	SB_T1_NORTH_SB_IN_B1,
	SB_T1_NORTH_SB_IN_B16,
	SB_T1_NORTH_SB_OUT_B1,
	SB_T1_NORTH_SB_OUT_B16,
	SB_T1_SOUTH_SB_IN_B1,
	SB_T1_SOUTH_SB_IN_B16,
	SB_T1_SOUTH_SB_OUT_B1,
	SB_T1_SOUTH_SB_OUT_B16,
	SB_T1_WEST_SB_IN_B1,
	SB_T1_WEST_SB_IN_B16,
	SB_T1_WEST_SB_OUT_B1,
	SB_T1_WEST_SB_OUT_B16,
	SB_T2_EAST_SB_IN_B1,
	SB_T2_EAST_SB_IN_B16,
	SB_T2_EAST_SB_OUT_B1,
	SB_T2_EAST_SB_OUT_B16,
	SB_T2_NORTH_SB_IN_B1,
	SB_T2_NORTH_SB_IN_B16,
	SB_T2_NORTH_SB_OUT_B1,
	SB_T2_NORTH_SB_OUT_B16,
	SB_T2_SOUTH_SB_IN_B1,
	SB_T2_SOUTH_SB_IN_B16,
	SB_T2_SOUTH_SB_OUT_B1,
	SB_T2_SOUTH_SB_OUT_B16,
	SB_T2_WEST_SB_IN_B1,
	SB_T2_WEST_SB_IN_B16,
	SB_T2_WEST_SB_OUT_B1,
	SB_T2_WEST_SB_OUT_B16,
	clk,
	clk_out,
	clk_pass_through,
	clk_pass_through_out_bot,
	config_config_addr,
	config_config_data,
	config_out_config_addr,
	config_out_config_data,
	config_out_read,
	config_out_write,
	config_read,
	config_write,
	hi,
	lo,
	read_config_data,
	read_config_data_in,
	reset,
	reset_out,
	stall,
	stall_out,
	tile_id
);
	input [0:0] SB_T0_EAST_SB_IN_B1;
	input [15:0] SB_T0_EAST_SB_IN_B16;
	output [0:0] SB_T0_EAST_SB_OUT_B1;
	output [15:0] SB_T0_EAST_SB_OUT_B16;
	input [0:0] SB_T0_NORTH_SB_IN_B1;
	input [15:0] SB_T0_NORTH_SB_IN_B16;
	output [0:0] SB_T0_NORTH_SB_OUT_B1;
	output [15:0] SB_T0_NORTH_SB_OUT_B16;
	input [0:0] SB_T0_SOUTH_SB_IN_B1;
	input [15:0] SB_T0_SOUTH_SB_IN_B16;
	output [0:0] SB_T0_SOUTH_SB_OUT_B1;
	output [15:0] SB_T0_SOUTH_SB_OUT_B16;
	input [0:0] SB_T0_WEST_SB_IN_B1;
	input [15:0] SB_T0_WEST_SB_IN_B16;
	output [0:0] SB_T0_WEST_SB_OUT_B1;
	output [15:0] SB_T0_WEST_SB_OUT_B16;
	input [0:0] SB_T1_EAST_SB_IN_B1;
	input [15:0] SB_T1_EAST_SB_IN_B16;
	output [0:0] SB_T1_EAST_SB_OUT_B1;
	output [15:0] SB_T1_EAST_SB_OUT_B16;
	input [0:0] SB_T1_NORTH_SB_IN_B1;
	input [15:0] SB_T1_NORTH_SB_IN_B16;
	output [0:0] SB_T1_NORTH_SB_OUT_B1;
	output [15:0] SB_T1_NORTH_SB_OUT_B16;
	input [0:0] SB_T1_SOUTH_SB_IN_B1;
	input [15:0] SB_T1_SOUTH_SB_IN_B16;
	output [0:0] SB_T1_SOUTH_SB_OUT_B1;
	output [15:0] SB_T1_SOUTH_SB_OUT_B16;
	input [0:0] SB_T1_WEST_SB_IN_B1;
	input [15:0] SB_T1_WEST_SB_IN_B16;
	output [0:0] SB_T1_WEST_SB_OUT_B1;
	output [15:0] SB_T1_WEST_SB_OUT_B16;
	input [0:0] SB_T2_EAST_SB_IN_B1;
	input [15:0] SB_T2_EAST_SB_IN_B16;
	output [0:0] SB_T2_EAST_SB_OUT_B1;
	output [15:0] SB_T2_EAST_SB_OUT_B16;
	input [0:0] SB_T2_NORTH_SB_IN_B1;
	input [15:0] SB_T2_NORTH_SB_IN_B16;
	output [0:0] SB_T2_NORTH_SB_OUT_B1;
	output [15:0] SB_T2_NORTH_SB_OUT_B16;
	input [0:0] SB_T2_SOUTH_SB_IN_B1;
	input [15:0] SB_T2_SOUTH_SB_IN_B16;
	output [0:0] SB_T2_SOUTH_SB_OUT_B1;
	output [15:0] SB_T2_SOUTH_SB_OUT_B16;
	input [0:0] SB_T2_WEST_SB_IN_B1;
	input [15:0] SB_T2_WEST_SB_IN_B16;
	output [0:0] SB_T2_WEST_SB_OUT_B1;
	output [15:0] SB_T2_WEST_SB_OUT_B16;
	input clk;
	output clk_out;
	input clk_pass_through;
	output clk_pass_through_out_bot;
	input [31:0] config_config_addr;
	input [31:0] config_config_data;
	output [31:0] config_out_config_addr;
	output [31:0] config_out_config_data;
	output [0:0] config_out_read;
	output [0:0] config_out_write;
	input [0:0] config_read;
	input [0:0] config_write;
	output [8:0] hi;
	output [7:0] lo;
	output [31:0] read_config_data;
	input [31:0] read_config_data_in;
	input reset;
	output reset_out;
	input [0:0] stall;
	output [0:0] stall_out;
	input [15:0] tile_id;
	wire [0:0] CB_bit0_O;
	wire [31:0] CB_bit0_read_config_data;
	wire [7:0] CB_bit0_config_config_addr_in;
	wire [0:0] CB_bit1_O;
	wire [31:0] CB_bit1_read_config_data;
	wire [7:0] CB_bit1_config_config_addr_in;
	wire [0:0] CB_bit2_O;
	wire [31:0] CB_bit2_read_config_data;
	wire [7:0] CB_bit2_config_config_addr_in;
	wire [15:0] CB_data0_O;
	wire [31:0] CB_data0_read_config_data;
	wire [7:0] CB_data0_config_config_addr_in;
	wire [15:0] CB_data1_O;
	wire [31:0] CB_data1_read_config_data;
	wire [7:0] CB_data1_config_config_addr_in;
	wire DECODE_FEATURE_0_O;
	wire DECODE_FEATURE_1_O;
	wire DECODE_FEATURE_2_O;
	wire DECODE_FEATURE_3_O;
	wire DECODE_FEATURE_4_O;
	wire DECODE_FEATURE_5_O;
	wire DECODE_FEATURE_6_O;
	wire DECODE_FEATURE_7_O;
	wire FEATURE_AND_0_out;
	wire FEATURE_AND_1_out;
	wire FEATURE_AND_2_out;
	wire FEATURE_AND_3_out;
	wire FEATURE_AND_4_out;
	wire FEATURE_AND_5_out;
	wire FEATURE_AND_6_out;
	wire FEATURE_AND_7_out;
	wire [15:0] PE_inst0_alu_res;
	wire [31:0] PE_inst0_read_config_data;
	wire [0:0] PE_inst0_res_p;
	wire [7:0] PE_inst0_config_config_addr_in;
	wire [15:0] SB_ID0_3TRACKS_B16_PE_SB_T0_EAST_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_PE_SB_T0_NORTH_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_PE_SB_T0_SOUTH_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_PE_SB_T0_WEST_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_PE_SB_T1_EAST_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_PE_SB_T1_NORTH_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_PE_SB_T1_SOUTH_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_PE_SB_T1_WEST_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_PE_SB_T2_EAST_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_PE_SB_T2_NORTH_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_PE_SB_T2_SOUTH_SB_OUT_B16;
	wire [15:0] SB_ID0_3TRACKS_B16_PE_SB_T2_WEST_SB_OUT_B16;
	wire [31:0] SB_ID0_3TRACKS_B16_PE_read_config_data;
	wire [7:0] SB_ID0_3TRACKS_B16_PE_config_config_addr_in;
	wire [0:0] SB_ID0_3TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1;
	wire [0:0] SB_ID0_3TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1;
	wire [31:0] SB_ID0_3TRACKS_B1_PE_read_config_data;
	wire [7:0] SB_ID0_3TRACKS_B1_PE_config_config_addr_in;
	wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T0_EAST_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T0_NORTH_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T0_SOUTH_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T0_WEST_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T1_EAST_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T1_NORTH_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T1_SOUTH_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T1_WEST_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T2_EAST_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T2_NORTH_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T2_SOUTH_SB_IN_B16_O;
	wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1_O;
	wire [15:0] WIRE_SB_T2_WEST_SB_IN_B16_O;
	wire and_inst0_out;
	wire and_inst1_out;
	wire [7:0] const_0_8_out;
	wire [8:0] const_511_9_out;
	wire coreir_eq_16_inst0_out;
	wire [31:0] read_config_data_or_inst0_out;
	wire [31:0] read_data_mux_O;
	wire [7:0] read_data_mux_S_in;
	wire [31:0] self_config_config_addr_out;
// diodes are put to prevent antenna violations on abutted pins
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T0 (.DIODE(tile_id[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T1 (.DIODE(tile_id[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T2 (.DIODE(tile_id[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T3 (.DIODE(tile_id[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T4 (.DIODE(tile_id[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T5 (.DIODE(tile_id[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T6 (.DIODE(tile_id[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T7 (.DIODE(tile_id[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T8 (.DIODE(tile_id[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T9 (.DIODE(tile_id[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T10 (.DIODE(tile_id[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T11 (.DIODE(tile_id[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T12 (.DIODE(tile_id[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T13 (.DIODE(tile_id[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T14 (.DIODE(tile_id[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_T15 (.DIODE(tile_id[15]));
// [start] input diodes
sky130_fd_sc_hd__diode_2 POHAN_DIODE_0 (.DIODE(SB_T0_EAST_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_1 (.DIODE(SB_T0_EAST_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_2 (.DIODE(SB_T0_EAST_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_3 (.DIODE(SB_T0_EAST_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_4 (.DIODE(SB_T0_EAST_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_5 (.DIODE(SB_T0_EAST_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_6 (.DIODE(SB_T0_EAST_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_7 (.DIODE(SB_T0_EAST_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_8 (.DIODE(SB_T0_EAST_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_9 (.DIODE(SB_T0_EAST_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_10 (.DIODE(SB_T0_EAST_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_11 (.DIODE(SB_T0_EAST_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_12 (.DIODE(SB_T0_EAST_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_13 (.DIODE(SB_T0_EAST_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_14 (.DIODE(SB_T0_EAST_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_15 (.DIODE(SB_T0_EAST_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_16 (.DIODE(SB_T0_EAST_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_17 (.DIODE(SB_T0_NORTH_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_18 (.DIODE(SB_T0_NORTH_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_19 (.DIODE(SB_T0_NORTH_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_20 (.DIODE(SB_T0_NORTH_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_21 (.DIODE(SB_T0_NORTH_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_22 (.DIODE(SB_T0_NORTH_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_23 (.DIODE(SB_T0_NORTH_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_24 (.DIODE(SB_T0_NORTH_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_25 (.DIODE(SB_T0_NORTH_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_26 (.DIODE(SB_T0_NORTH_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_27 (.DIODE(SB_T0_NORTH_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_28 (.DIODE(SB_T0_NORTH_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_29 (.DIODE(SB_T0_NORTH_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_30 (.DIODE(SB_T0_NORTH_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_31 (.DIODE(SB_T0_NORTH_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_32 (.DIODE(SB_T0_NORTH_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_33 (.DIODE(SB_T0_NORTH_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_34 (.DIODE(SB_T0_SOUTH_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_35 (.DIODE(SB_T0_SOUTH_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_36 (.DIODE(SB_T0_SOUTH_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_37 (.DIODE(SB_T0_SOUTH_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_38 (.DIODE(SB_T0_SOUTH_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_39 (.DIODE(SB_T0_SOUTH_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_40 (.DIODE(SB_T0_SOUTH_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_41 (.DIODE(SB_T0_SOUTH_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_42 (.DIODE(SB_T0_SOUTH_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_43 (.DIODE(SB_T0_SOUTH_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_44 (.DIODE(SB_T0_SOUTH_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_45 (.DIODE(SB_T0_SOUTH_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_46 (.DIODE(SB_T0_SOUTH_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_47 (.DIODE(SB_T0_SOUTH_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_48 (.DIODE(SB_T0_SOUTH_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_49 (.DIODE(SB_T0_SOUTH_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_50 (.DIODE(SB_T0_SOUTH_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_51 (.DIODE(SB_T0_WEST_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_52 (.DIODE(SB_T0_WEST_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_53 (.DIODE(SB_T0_WEST_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_54 (.DIODE(SB_T0_WEST_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_55 (.DIODE(SB_T0_WEST_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_56 (.DIODE(SB_T0_WEST_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_57 (.DIODE(SB_T0_WEST_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_58 (.DIODE(SB_T0_WEST_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_59 (.DIODE(SB_T0_WEST_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_60 (.DIODE(SB_T0_WEST_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_61 (.DIODE(SB_T0_WEST_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_62 (.DIODE(SB_T0_WEST_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_63 (.DIODE(SB_T0_WEST_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_64 (.DIODE(SB_T0_WEST_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_65 (.DIODE(SB_T0_WEST_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_66 (.DIODE(SB_T0_WEST_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_67 (.DIODE(SB_T0_WEST_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_68 (.DIODE(SB_T1_EAST_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_69 (.DIODE(SB_T1_EAST_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_70 (.DIODE(SB_T1_EAST_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_71 (.DIODE(SB_T1_EAST_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_72 (.DIODE(SB_T1_EAST_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_73 (.DIODE(SB_T1_EAST_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_74 (.DIODE(SB_T1_EAST_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_75 (.DIODE(SB_T1_EAST_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_76 (.DIODE(SB_T1_EAST_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_77 (.DIODE(SB_T1_EAST_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_78 (.DIODE(SB_T1_EAST_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_79 (.DIODE(SB_T1_EAST_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_80 (.DIODE(SB_T1_EAST_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_81 (.DIODE(SB_T1_EAST_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_82 (.DIODE(SB_T1_EAST_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_83 (.DIODE(SB_T1_EAST_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_84 (.DIODE(SB_T1_EAST_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_85 (.DIODE(SB_T1_NORTH_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_86 (.DIODE(SB_T1_NORTH_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_87 (.DIODE(SB_T1_NORTH_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_88 (.DIODE(SB_T1_NORTH_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_89 (.DIODE(SB_T1_NORTH_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_90 (.DIODE(SB_T1_NORTH_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_91 (.DIODE(SB_T1_NORTH_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_92 (.DIODE(SB_T1_NORTH_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_93 (.DIODE(SB_T1_NORTH_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_94 (.DIODE(SB_T1_NORTH_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_95 (.DIODE(SB_T1_NORTH_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_96 (.DIODE(SB_T1_NORTH_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_97 (.DIODE(SB_T1_NORTH_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_98 (.DIODE(SB_T1_NORTH_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_99 (.DIODE(SB_T1_NORTH_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_100 (.DIODE(SB_T1_NORTH_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_101 (.DIODE(SB_T1_NORTH_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_102 (.DIODE(SB_T1_SOUTH_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_103 (.DIODE(SB_T1_SOUTH_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_104 (.DIODE(SB_T1_SOUTH_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_105 (.DIODE(SB_T1_SOUTH_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_106 (.DIODE(SB_T1_SOUTH_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_107 (.DIODE(SB_T1_SOUTH_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_108 (.DIODE(SB_T1_SOUTH_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_109 (.DIODE(SB_T1_SOUTH_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_110 (.DIODE(SB_T1_SOUTH_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_111 (.DIODE(SB_T1_SOUTH_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_112 (.DIODE(SB_T1_SOUTH_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_113 (.DIODE(SB_T1_SOUTH_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_114 (.DIODE(SB_T1_SOUTH_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_115 (.DIODE(SB_T1_SOUTH_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_116 (.DIODE(SB_T1_SOUTH_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_117 (.DIODE(SB_T1_SOUTH_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_118 (.DIODE(SB_T1_SOUTH_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_119 (.DIODE(SB_T1_WEST_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_120 (.DIODE(SB_T1_WEST_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_121 (.DIODE(SB_T1_WEST_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_122 (.DIODE(SB_T1_WEST_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_123 (.DIODE(SB_T1_WEST_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_124 (.DIODE(SB_T1_WEST_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_125 (.DIODE(SB_T1_WEST_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_126 (.DIODE(SB_T1_WEST_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_127 (.DIODE(SB_T1_WEST_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_128 (.DIODE(SB_T1_WEST_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_129 (.DIODE(SB_T1_WEST_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_130 (.DIODE(SB_T1_WEST_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_131 (.DIODE(SB_T1_WEST_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_132 (.DIODE(SB_T1_WEST_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_133 (.DIODE(SB_T1_WEST_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_134 (.DIODE(SB_T1_WEST_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_135 (.DIODE(SB_T1_WEST_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_136 (.DIODE(SB_T2_EAST_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_137 (.DIODE(SB_T2_EAST_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_138 (.DIODE(SB_T2_EAST_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_139 (.DIODE(SB_T2_EAST_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_140 (.DIODE(SB_T2_EAST_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_141 (.DIODE(SB_T2_EAST_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_142 (.DIODE(SB_T2_EAST_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_143 (.DIODE(SB_T2_EAST_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_144 (.DIODE(SB_T2_EAST_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_145 (.DIODE(SB_T2_EAST_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_146 (.DIODE(SB_T2_EAST_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_147 (.DIODE(SB_T2_EAST_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_148 (.DIODE(SB_T2_EAST_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_149 (.DIODE(SB_T2_EAST_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_150 (.DIODE(SB_T2_EAST_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_151 (.DIODE(SB_T2_EAST_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_152 (.DIODE(SB_T2_EAST_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_153 (.DIODE(SB_T2_NORTH_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_154 (.DIODE(SB_T2_NORTH_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_155 (.DIODE(SB_T2_NORTH_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_156 (.DIODE(SB_T2_NORTH_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_157 (.DIODE(SB_T2_NORTH_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_158 (.DIODE(SB_T2_NORTH_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_159 (.DIODE(SB_T2_NORTH_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_160 (.DIODE(SB_T2_NORTH_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_161 (.DIODE(SB_T2_NORTH_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_162 (.DIODE(SB_T2_NORTH_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_163 (.DIODE(SB_T2_NORTH_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_164 (.DIODE(SB_T2_NORTH_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_165 (.DIODE(SB_T2_NORTH_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_166 (.DIODE(SB_T2_NORTH_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_167 (.DIODE(SB_T2_NORTH_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_168 (.DIODE(SB_T2_NORTH_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_169 (.DIODE(SB_T2_NORTH_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_170 (.DIODE(SB_T2_SOUTH_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_171 (.DIODE(SB_T2_SOUTH_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_172 (.DIODE(SB_T2_SOUTH_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_173 (.DIODE(SB_T2_SOUTH_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_174 (.DIODE(SB_T2_SOUTH_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_175 (.DIODE(SB_T2_SOUTH_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_176 (.DIODE(SB_T2_SOUTH_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_177 (.DIODE(SB_T2_SOUTH_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_178 (.DIODE(SB_T2_SOUTH_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_179 (.DIODE(SB_T2_SOUTH_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_180 (.DIODE(SB_T2_SOUTH_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_181 (.DIODE(SB_T2_SOUTH_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_182 (.DIODE(SB_T2_SOUTH_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_183 (.DIODE(SB_T2_SOUTH_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_184 (.DIODE(SB_T2_SOUTH_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_185 (.DIODE(SB_T2_SOUTH_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_186 (.DIODE(SB_T2_SOUTH_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_187 (.DIODE(SB_T2_WEST_SB_IN_B1[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_188 (.DIODE(SB_T2_WEST_SB_IN_B16[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_189 (.DIODE(SB_T2_WEST_SB_IN_B16[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_190 (.DIODE(SB_T2_WEST_SB_IN_B16[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_191 (.DIODE(SB_T2_WEST_SB_IN_B16[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_192 (.DIODE(SB_T2_WEST_SB_IN_B16[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_193 (.DIODE(SB_T2_WEST_SB_IN_B16[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_194 (.DIODE(SB_T2_WEST_SB_IN_B16[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_195 (.DIODE(SB_T2_WEST_SB_IN_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_196 (.DIODE(SB_T2_WEST_SB_IN_B16[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_197 (.DIODE(SB_T2_WEST_SB_IN_B16[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_198 (.DIODE(SB_T2_WEST_SB_IN_B16[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_199 (.DIODE(SB_T2_WEST_SB_IN_B16[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_200 (.DIODE(SB_T2_WEST_SB_IN_B16[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_201 (.DIODE(SB_T2_WEST_SB_IN_B16[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_202 (.DIODE(SB_T2_WEST_SB_IN_B16[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_203 (.DIODE(SB_T2_WEST_SB_IN_B16[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_204 (.DIODE(clk));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_205 (.DIODE(clk_pass_through));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_206 (.DIODE(config_config_addr[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_207 (.DIODE(config_config_addr[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_208 (.DIODE(config_config_addr[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_209 (.DIODE(config_config_addr[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_210 (.DIODE(config_config_addr[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_211 (.DIODE(config_config_addr[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_212 (.DIODE(config_config_addr[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_213 (.DIODE(config_config_addr[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_214 (.DIODE(config_config_addr[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_215 (.DIODE(config_config_addr[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_216 (.DIODE(config_config_addr[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_217 (.DIODE(config_config_addr[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_218 (.DIODE(config_config_addr[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_219 (.DIODE(config_config_addr[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_220 (.DIODE(config_config_addr[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_221 (.DIODE(config_config_addr[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_222 (.DIODE(config_config_addr[16]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_223 (.DIODE(config_config_addr[17]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_224 (.DIODE(config_config_addr[18]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_225 (.DIODE(config_config_addr[19]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_226 (.DIODE(config_config_addr[20]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_227 (.DIODE(config_config_addr[21]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_228 (.DIODE(config_config_addr[22]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_229 (.DIODE(config_config_addr[23]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_230 (.DIODE(config_config_addr[24]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_231 (.DIODE(config_config_addr[25]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_232 (.DIODE(config_config_addr[26]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_233 (.DIODE(config_config_addr[27]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_234 (.DIODE(config_config_addr[28]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_235 (.DIODE(config_config_addr[29]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_236 (.DIODE(config_config_addr[30]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_237 (.DIODE(config_config_addr[31]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_238 (.DIODE(config_config_data[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_239 (.DIODE(config_config_data[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_240 (.DIODE(config_config_data[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_241 (.DIODE(config_config_data[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_242 (.DIODE(config_config_data[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_243 (.DIODE(config_config_data[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_244 (.DIODE(config_config_data[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_245 (.DIODE(config_config_data[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_246 (.DIODE(config_config_data[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_247 (.DIODE(config_config_data[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_248 (.DIODE(config_config_data[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_249 (.DIODE(config_config_data[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_250 (.DIODE(config_config_data[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_251 (.DIODE(config_config_data[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_252 (.DIODE(config_config_data[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_253 (.DIODE(config_config_data[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_254 (.DIODE(config_config_data[16]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_255 (.DIODE(config_config_data[17]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_256 (.DIODE(config_config_data[18]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_257 (.DIODE(config_config_data[19]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_258 (.DIODE(config_config_data[20]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_259 (.DIODE(config_config_data[21]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_260 (.DIODE(config_config_data[22]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_261 (.DIODE(config_config_data[23]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_262 (.DIODE(config_config_data[24]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_263 (.DIODE(config_config_data[25]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_264 (.DIODE(config_config_data[26]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_265 (.DIODE(config_config_data[27]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_266 (.DIODE(config_config_data[28]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_267 (.DIODE(config_config_data[29]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_268 (.DIODE(config_config_data[30]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_269 (.DIODE(config_config_data[31]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_270 (.DIODE(config_read[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_271 (.DIODE(config_write[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_272 (.DIODE(read_config_data_in[0]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_273 (.DIODE(read_config_data_in[1]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_274 (.DIODE(read_config_data_in[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_275 (.DIODE(read_config_data_in[3]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_276 (.DIODE(read_config_data_in[4]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_277 (.DIODE(read_config_data_in[5]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_278 (.DIODE(read_config_data_in[6]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_279 (.DIODE(read_config_data_in[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_280 (.DIODE(read_config_data_in[8]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_281 (.DIODE(read_config_data_in[9]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_282 (.DIODE(read_config_data_in[10]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_283 (.DIODE(read_config_data_in[11]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_284 (.DIODE(read_config_data_in[12]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_285 (.DIODE(read_config_data_in[13]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_286 (.DIODE(read_config_data_in[14]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_287 (.DIODE(read_config_data_in[15]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_288 (.DIODE(read_config_data_in[16]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_289 (.DIODE(read_config_data_in[17]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_290 (.DIODE(read_config_data_in[18]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_291 (.DIODE(read_config_data_in[19]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_292 (.DIODE(read_config_data_in[20]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_293 (.DIODE(read_config_data_in[21]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_294 (.DIODE(read_config_data_in[22]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_295 (.DIODE(read_config_data_in[23]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_296 (.DIODE(read_config_data_in[24]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_297 (.DIODE(read_config_data_in[25]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_298 (.DIODE(read_config_data_in[26]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_299 (.DIODE(read_config_data_in[27]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_300 (.DIODE(read_config_data_in[28]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_301 (.DIODE(read_config_data_in[29]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_302 (.DIODE(read_config_data_in[30]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_303 (.DIODE(read_config_data_in[31]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_304 (.DIODE(reset));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_305 (.DIODE(stall[0]));
// [end] input diodes

// [start] output diodes
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_306 (.DIODE(SB_T0_EAST_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_307 (.DIODE(SB_T0_EAST_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_308 (.DIODE(SB_T0_EAST_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_309 (.DIODE(SB_T0_EAST_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_310 (.DIODE(SB_T0_EAST_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_311 (.DIODE(SB_T0_EAST_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_312 (.DIODE(SB_T0_EAST_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_313 (.DIODE(SB_T0_EAST_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_314 (.DIODE(SB_T0_EAST_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_315 (.DIODE(SB_T0_EAST_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_316 (.DIODE(SB_T0_EAST_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_317 (.DIODE(SB_T0_EAST_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_318 (.DIODE(SB_T0_EAST_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_319 (.DIODE(SB_T0_EAST_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_320 (.DIODE(SB_T0_EAST_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_321 (.DIODE(SB_T0_EAST_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_322 (.DIODE(SB_T0_EAST_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_323 (.DIODE(SB_T0_NORTH_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_324 (.DIODE(SB_T0_NORTH_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_325 (.DIODE(SB_T0_NORTH_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_326 (.DIODE(SB_T0_NORTH_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_327 (.DIODE(SB_T0_NORTH_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_328 (.DIODE(SB_T0_NORTH_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_329 (.DIODE(SB_T0_NORTH_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_330 (.DIODE(SB_T0_NORTH_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_331 (.DIODE(SB_T0_NORTH_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_332 (.DIODE(SB_T0_NORTH_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_333 (.DIODE(SB_T0_NORTH_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_334 (.DIODE(SB_T0_NORTH_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_335 (.DIODE(SB_T0_NORTH_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_336 (.DIODE(SB_T0_NORTH_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_337 (.DIODE(SB_T0_NORTH_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_338 (.DIODE(SB_T0_NORTH_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_339 (.DIODE(SB_T0_NORTH_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_340 (.DIODE(SB_T0_SOUTH_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_341 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_342 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_343 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_344 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_345 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_346 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_347 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_348 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_349 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_350 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_351 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_352 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_353 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_354 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_355 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_356 (.DIODE(SB_T0_SOUTH_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_357 (.DIODE(SB_T0_WEST_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_358 (.DIODE(SB_T0_WEST_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_359 (.DIODE(SB_T0_WEST_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_360 (.DIODE(SB_T0_WEST_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_361 (.DIODE(SB_T0_WEST_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_362 (.DIODE(SB_T0_WEST_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_363 (.DIODE(SB_T0_WEST_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_364 (.DIODE(SB_T0_WEST_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_365 (.DIODE(SB_T0_WEST_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_366 (.DIODE(SB_T0_WEST_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_367 (.DIODE(SB_T0_WEST_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_368 (.DIODE(SB_T0_WEST_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_369 (.DIODE(SB_T0_WEST_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_370 (.DIODE(SB_T0_WEST_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_371 (.DIODE(SB_T0_WEST_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_372 (.DIODE(SB_T0_WEST_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_373 (.DIODE(SB_T0_WEST_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_374 (.DIODE(SB_T1_EAST_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_375 (.DIODE(SB_T1_EAST_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_376 (.DIODE(SB_T1_EAST_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_377 (.DIODE(SB_T1_EAST_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_378 (.DIODE(SB_T1_EAST_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_379 (.DIODE(SB_T1_EAST_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_380 (.DIODE(SB_T1_EAST_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_381 (.DIODE(SB_T1_EAST_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_382 (.DIODE(SB_T1_EAST_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_383 (.DIODE(SB_T1_EAST_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_384 (.DIODE(SB_T1_EAST_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_385 (.DIODE(SB_T1_EAST_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_386 (.DIODE(SB_T1_EAST_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_387 (.DIODE(SB_T1_EAST_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_388 (.DIODE(SB_T1_EAST_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_389 (.DIODE(SB_T1_EAST_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_390 (.DIODE(SB_T1_EAST_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_391 (.DIODE(SB_T1_NORTH_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_392 (.DIODE(SB_T1_NORTH_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_393 (.DIODE(SB_T1_NORTH_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_394 (.DIODE(SB_T1_NORTH_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_395 (.DIODE(SB_T1_NORTH_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_396 (.DIODE(SB_T1_NORTH_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_397 (.DIODE(SB_T1_NORTH_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_398 (.DIODE(SB_T1_NORTH_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_399 (.DIODE(SB_T1_NORTH_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_400 (.DIODE(SB_T1_NORTH_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_401 (.DIODE(SB_T1_NORTH_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_402 (.DIODE(SB_T1_NORTH_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_403 (.DIODE(SB_T1_NORTH_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_404 (.DIODE(SB_T1_NORTH_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_405 (.DIODE(SB_T1_NORTH_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_406 (.DIODE(SB_T1_NORTH_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_407 (.DIODE(SB_T1_NORTH_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_408 (.DIODE(SB_T1_SOUTH_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_409 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_410 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_411 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_412 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_413 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_414 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_415 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_416 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_417 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_418 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_419 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_420 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_421 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_422 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_423 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_424 (.DIODE(SB_T1_SOUTH_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_425 (.DIODE(SB_T1_WEST_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_426 (.DIODE(SB_T1_WEST_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_427 (.DIODE(SB_T1_WEST_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_428 (.DIODE(SB_T1_WEST_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_429 (.DIODE(SB_T1_WEST_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_430 (.DIODE(SB_T1_WEST_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_431 (.DIODE(SB_T1_WEST_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_432 (.DIODE(SB_T1_WEST_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_433 (.DIODE(SB_T1_WEST_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_434 (.DIODE(SB_T1_WEST_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_435 (.DIODE(SB_T1_WEST_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_436 (.DIODE(SB_T1_WEST_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_437 (.DIODE(SB_T1_WEST_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_438 (.DIODE(SB_T1_WEST_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_439 (.DIODE(SB_T1_WEST_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_440 (.DIODE(SB_T1_WEST_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_441 (.DIODE(SB_T1_WEST_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_442 (.DIODE(SB_T2_EAST_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_443 (.DIODE(SB_T2_EAST_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_444 (.DIODE(SB_T2_EAST_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_445 (.DIODE(SB_T2_EAST_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_446 (.DIODE(SB_T2_EAST_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_447 (.DIODE(SB_T2_EAST_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_448 (.DIODE(SB_T2_EAST_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_449 (.DIODE(SB_T2_EAST_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_450 (.DIODE(SB_T2_EAST_SB_OUT_B16[7]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_451 (.DIODE(SB_T2_EAST_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_452 (.DIODE(SB_T2_EAST_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_453 (.DIODE(SB_T2_EAST_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_454 (.DIODE(SB_T2_EAST_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_455 (.DIODE(SB_T2_EAST_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_456 (.DIODE(SB_T2_EAST_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_457 (.DIODE(SB_T2_EAST_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_458 (.DIODE(SB_T2_EAST_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_459 (.DIODE(SB_T2_NORTH_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_460 (.DIODE(SB_T2_NORTH_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_461 (.DIODE(SB_T2_NORTH_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_462 (.DIODE(SB_T2_NORTH_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_463 (.DIODE(SB_T2_NORTH_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_464 (.DIODE(SB_T2_NORTH_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_465 (.DIODE(SB_T2_NORTH_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_466 (.DIODE(SB_T2_NORTH_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_467 (.DIODE(SB_T2_NORTH_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_468 (.DIODE(SB_T2_NORTH_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_469 (.DIODE(SB_T2_NORTH_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_470 (.DIODE(SB_T2_NORTH_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_471 (.DIODE(SB_T2_NORTH_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_472 (.DIODE(SB_T2_NORTH_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_473 (.DIODE(SB_T2_NORTH_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_474 (.DIODE(SB_T2_NORTH_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_475 (.DIODE(SB_T2_NORTH_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_476 (.DIODE(SB_T2_SOUTH_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_477 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_478 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_479 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_480 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_481 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_482 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_483 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_484 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_485 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_486 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_487 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_488 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_489 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_490 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_491 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_492 (.DIODE(SB_T2_SOUTH_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_493 (.DIODE(SB_T2_WEST_SB_OUT_B1[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_494 (.DIODE(SB_T2_WEST_SB_OUT_B16[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_495 (.DIODE(SB_T2_WEST_SB_OUT_B16[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_496 (.DIODE(SB_T2_WEST_SB_OUT_B16[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_497 (.DIODE(SB_T2_WEST_SB_OUT_B16[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_498 (.DIODE(SB_T2_WEST_SB_OUT_B16[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_499 (.DIODE(SB_T2_WEST_SB_OUT_B16[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_500 (.DIODE(SB_T2_WEST_SB_OUT_B16[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_501 (.DIODE(SB_T2_WEST_SB_OUT_B16[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_502 (.DIODE(SB_T2_WEST_SB_OUT_B16[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_503 (.DIODE(SB_T2_WEST_SB_OUT_B16[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_504 (.DIODE(SB_T2_WEST_SB_OUT_B16[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_505 (.DIODE(SB_T2_WEST_SB_OUT_B16[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_506 (.DIODE(SB_T2_WEST_SB_OUT_B16[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_507 (.DIODE(SB_T2_WEST_SB_OUT_B16[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_508 (.DIODE(SB_T2_WEST_SB_OUT_B16[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_509 (.DIODE(SB_T2_WEST_SB_OUT_B16[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_510 (.DIODE(clk_out));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_511 (.DIODE(clk_pass_through_out_bot));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_512 (.DIODE(config_out_config_addr[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_513 (.DIODE(config_out_config_addr[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_514 (.DIODE(config_out_config_addr[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_515 (.DIODE(config_out_config_addr[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_516 (.DIODE(config_out_config_addr[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_517 (.DIODE(config_out_config_addr[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_518 (.DIODE(config_out_config_addr[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_519 (.DIODE(config_out_config_addr[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_520 (.DIODE(config_out_config_addr[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_521 (.DIODE(config_out_config_addr[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_522 (.DIODE(config_out_config_addr[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_523 (.DIODE(config_out_config_addr[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_524 (.DIODE(config_out_config_addr[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_525 (.DIODE(config_out_config_addr[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_526 (.DIODE(config_out_config_addr[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_527 (.DIODE(config_out_config_addr[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_528 (.DIODE(config_out_config_addr[16]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_529 (.DIODE(config_out_config_addr[17]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_530 (.DIODE(config_out_config_addr[18]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_531 (.DIODE(config_out_config_addr[19]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_532 (.DIODE(config_out_config_addr[20]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_533 (.DIODE(config_out_config_addr[21]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_534 (.DIODE(config_out_config_addr[22]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_535 (.DIODE(config_out_config_addr[23]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_536 (.DIODE(config_out_config_addr[24]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_537 (.DIODE(config_out_config_addr[25]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_538 (.DIODE(config_out_config_addr[26]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_539 (.DIODE(config_out_config_addr[27]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_540 (.DIODE(config_out_config_addr[28]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_541 (.DIODE(config_out_config_addr[29]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_542 (.DIODE(config_out_config_addr[30]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_543 (.DIODE(config_out_config_addr[31]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_544 (.DIODE(config_out_config_data[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_545 (.DIODE(config_out_config_data[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_546 (.DIODE(config_out_config_data[2]));
sky130_fd_sc_hd__diode_2 POHAN_DIODE_547 (.DIODE(config_out_config_data[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_548 (.DIODE(config_out_config_data[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_549 (.DIODE(config_out_config_data[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_550 (.DIODE(config_out_config_data[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_551 (.DIODE(config_out_config_data[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_552 (.DIODE(config_out_config_data[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_553 (.DIODE(config_out_config_data[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_554 (.DIODE(config_out_config_data[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_555 (.DIODE(config_out_config_data[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_556 (.DIODE(config_out_config_data[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_557 (.DIODE(config_out_config_data[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_558 (.DIODE(config_out_config_data[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_559 (.DIODE(config_out_config_data[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_560 (.DIODE(config_out_config_data[16]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_561 (.DIODE(config_out_config_data[17]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_562 (.DIODE(config_out_config_data[18]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_563 (.DIODE(config_out_config_data[19]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_564 (.DIODE(config_out_config_data[20]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_565 (.DIODE(config_out_config_data[21]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_566 (.DIODE(config_out_config_data[22]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_567 (.DIODE(config_out_config_data[23]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_568 (.DIODE(config_out_config_data[24]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_569 (.DIODE(config_out_config_data[25]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_570 (.DIODE(config_out_config_data[26]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_571 (.DIODE(config_out_config_data[27]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_572 (.DIODE(config_out_config_data[28]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_573 (.DIODE(config_out_config_data[29]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_574 (.DIODE(config_out_config_data[30]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_575 (.DIODE(config_out_config_data[31]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_576 (.DIODE(config_out_read[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_577 (.DIODE(config_out_write[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_578 (.DIODE(read_config_data[0]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_579 (.DIODE(read_config_data[1]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_580 (.DIODE(read_config_data[2]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_581 (.DIODE(read_config_data[3]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_582 (.DIODE(read_config_data[4]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_583 (.DIODE(read_config_data[5]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_584 (.DIODE(read_config_data[6]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_585 (.DIODE(read_config_data[7]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_586 (.DIODE(read_config_data[8]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_587 (.DIODE(read_config_data[9]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_588 (.DIODE(read_config_data[10]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_589 (.DIODE(read_config_data[11]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_590 (.DIODE(read_config_data[12]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_591 (.DIODE(read_config_data[13]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_592 (.DIODE(read_config_data[14]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_593 (.DIODE(read_config_data[15]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_594 (.DIODE(read_config_data[16]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_595 (.DIODE(read_config_data[17]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_596 (.DIODE(read_config_data[18]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_597 (.DIODE(read_config_data[19]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_598 (.DIODE(read_config_data[20]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_599 (.DIODE(read_config_data[21]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_600 (.DIODE(read_config_data[22]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_601 (.DIODE(read_config_data[23]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_602 (.DIODE(read_config_data[24]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_603 (.DIODE(read_config_data[25]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_604 (.DIODE(read_config_data[26]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_605 (.DIODE(read_config_data[27]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_606 (.DIODE(read_config_data[28]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_607 (.DIODE(read_config_data[29]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_608 (.DIODE(read_config_data[30]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_609 (.DIODE(read_config_data[31]));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_610 (.DIODE(reset_out));
// sky130_fd_sc_hd__diode_2 POHAN_DIODE_611 (.DIODE(stall_out[0]));
// [end] output diodes
	CB_bit0 CB_bit0(
		.I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
		.I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
		.I_10(WIRE_SB_T2_EAST_SB_IN_B1_O),
		.I_11(WIRE_SB_T2_WEST_SB_IN_B1_O),
		.I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
		.I_3(WIRE_SB_T0_WEST_SB_IN_B1_O),
		.I_4(WIRE_SB_T1_NORTH_SB_IN_B1_O),
		.I_5(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
		.I_6(WIRE_SB_T1_EAST_SB_IN_B1_O),
		.I_7(WIRE_SB_T1_WEST_SB_IN_B1_O),
		.I_8(WIRE_SB_T2_NORTH_SB_IN_B1_O),
		.I_9(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
		.O(CB_bit0_O),
		.clk(clk),
		.config_config_addr(CB_bit0_config_config_addr_in),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_1_out),
		.read_config_data(CB_bit0_read_config_data),
		.reset(reset)
	);
	mantle_wire__typeBitIn8 CB_bit0_config_config_addr(
		.in(CB_bit0_config_config_addr_in),
		.out(self_config_config_addr_out[31:24])
	);
	CB_bit1 CB_bit1(
		.I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
		.I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
		.I_10(WIRE_SB_T2_EAST_SB_IN_B1_O),
		.I_11(WIRE_SB_T2_WEST_SB_IN_B1_O),
		.I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
		.I_3(WIRE_SB_T0_WEST_SB_IN_B1_O),
		.I_4(WIRE_SB_T1_NORTH_SB_IN_B1_O),
		.I_5(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
		.I_6(WIRE_SB_T1_EAST_SB_IN_B1_O),
		.I_7(WIRE_SB_T1_WEST_SB_IN_B1_O),
		.I_8(WIRE_SB_T2_NORTH_SB_IN_B1_O),
		.I_9(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
		.O(CB_bit1_O),
		.clk(clk),
		.config_config_addr(CB_bit1_config_config_addr_in),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_2_out),
		.read_config_data(CB_bit1_read_config_data),
		.reset(reset)
	);
	mantle_wire__typeBitIn8 CB_bit1_config_config_addr(
		.in(CB_bit1_config_config_addr_in),
		.out(self_config_config_addr_out[31:24])
	);
	CB_bit2 CB_bit2(
		.I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
		.I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
		.I_10(WIRE_SB_T2_EAST_SB_IN_B1_O),
		.I_11(WIRE_SB_T2_WEST_SB_IN_B1_O),
		.I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
		.I_3(WIRE_SB_T0_WEST_SB_IN_B1_O),
		.I_4(WIRE_SB_T1_NORTH_SB_IN_B1_O),
		.I_5(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
		.I_6(WIRE_SB_T1_EAST_SB_IN_B1_O),
		.I_7(WIRE_SB_T1_WEST_SB_IN_B1_O),
		.I_8(WIRE_SB_T2_NORTH_SB_IN_B1_O),
		.I_9(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
		.O(CB_bit2_O),
		.clk(clk),
		.config_config_addr(CB_bit2_config_config_addr_in),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_3_out),
		.read_config_data(CB_bit2_read_config_data),
		.reset(reset)
	);
	mantle_wire__typeBitIn8 CB_bit2_config_config_addr(
		.in(CB_bit2_config_config_addr_in),
		.out(self_config_config_addr_out[31:24])
	);
	CB_data0 CB_data0(
		.I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
		.I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
		.I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
		.I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
		.I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
		.I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
		.I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
		.I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
		.I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
		.I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
		.I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
		.I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
		.O(CB_data0_O),
		.clk(clk),
		.config_config_addr(CB_data0_config_config_addr_in),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_4_out),
		.read_config_data(CB_data0_read_config_data),
		.reset(reset)
	);
	mantle_wire__typeBitIn8 CB_data0_config_config_addr(
		.in(CB_data0_config_config_addr_in),
		.out(self_config_config_addr_out[31:24])
	);
	CB_data1 CB_data1(
		.I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
		.I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
		.I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
		.I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
		.I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
		.I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
		.I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
		.I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
		.I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
		.I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
		.I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
		.I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
		.O(CB_data1_O),
		.clk(clk),
		.config_config_addr(CB_data1_config_config_addr_in),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_5_out),
		.read_config_data(CB_data1_read_config_data),
		.reset(reset)
	);
	mantle_wire__typeBitIn8 CB_data1_config_config_addr(
		.in(CB_data1_config_config_addr_in),
		.out(self_config_config_addr_out[31:24])
	);
	Decode08 DECODE_FEATURE_0(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_0_O)
	);
	Decode18 DECODE_FEATURE_1(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_1_O)
	);
	Decode28 DECODE_FEATURE_2(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_2_O)
	);
	Decode38 DECODE_FEATURE_3(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_3_O)
	);
	Decode48 DECODE_FEATURE_4(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_4_O)
	);
	Decode58 DECODE_FEATURE_5(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_5_O)
	);
	Decode68 DECODE_FEATURE_6(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_6_O)
	);
	Decode78 DECODE_FEATURE_7(
		.I(self_config_config_addr_out[23:16]),
		.O(DECODE_FEATURE_7_O)
	);
	corebit_and FEATURE_AND_0(
		.in0(DECODE_FEATURE_0_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_0_out)
	);
	corebit_and FEATURE_AND_1(
		.in0(DECODE_FEATURE_1_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_1_out)
	);
	corebit_and FEATURE_AND_2(
		.in0(DECODE_FEATURE_2_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_2_out)
	);
	corebit_and FEATURE_AND_3(
		.in0(DECODE_FEATURE_3_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_3_out)
	);
	corebit_and FEATURE_AND_4(
		.in0(DECODE_FEATURE_4_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_4_out)
	);
	corebit_and FEATURE_AND_5(
		.in0(DECODE_FEATURE_5_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_5_out)
	);
	corebit_and FEATURE_AND_6(
		.in0(DECODE_FEATURE_6_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_6_out)
	);
	corebit_and FEATURE_AND_7(
		.in0(DECODE_FEATURE_7_O),
		.in1(and_inst1_out),
		.out(FEATURE_AND_7_out)
	);
	PE_unq1 PE_inst0(
		.alu_res(PE_inst0_alu_res),
		.bit0(CB_bit0_O),
		.bit1(CB_bit1_O),
		.bit2(CB_bit2_O),
		.clk(clk),
		.config_config_addr(PE_inst0_config_config_addr_in),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_0_out),
		.data0(CB_data0_O),
		.data1(CB_data1_O),
		.read_config_data(PE_inst0_read_config_data),
		.res_p(PE_inst0_res_p),
		.reset(reset),
		.stall(stall)
	);
	mantle_wire__typeBitIn8 PE_inst0_config_config_addr(
		.in(PE_inst0_config_config_addr_in),
		.out(self_config_config_addr_out[31:24])
	);
	SB_ID0_3TRACKS_B16_PE SB_ID0_3TRACKS_B16_PE(
		.SB_T0_EAST_SB_IN_B16(SB_T0_EAST_SB_IN_B16),
		.SB_T0_EAST_SB_OUT_B16(SB_ID0_3TRACKS_B16_PE_SB_T0_EAST_SB_OUT_B16),
		.SB_T0_NORTH_SB_IN_B16(SB_T0_NORTH_SB_IN_B16),
		.SB_T0_NORTH_SB_OUT_B16(SB_ID0_3TRACKS_B16_PE_SB_T0_NORTH_SB_OUT_B16),
		.SB_T0_SOUTH_SB_IN_B16(SB_T0_SOUTH_SB_IN_B16),
		.SB_T0_SOUTH_SB_OUT_B16(SB_ID0_3TRACKS_B16_PE_SB_T0_SOUTH_SB_OUT_B16),
		.SB_T0_WEST_SB_IN_B16(SB_T0_WEST_SB_IN_B16),
		.SB_T0_WEST_SB_OUT_B16(SB_ID0_3TRACKS_B16_PE_SB_T0_WEST_SB_OUT_B16),
		.SB_T1_EAST_SB_IN_B16(SB_T1_EAST_SB_IN_B16),
		.SB_T1_EAST_SB_OUT_B16(SB_ID0_3TRACKS_B16_PE_SB_T1_EAST_SB_OUT_B16),
		.SB_T1_NORTH_SB_IN_B16(SB_T1_NORTH_SB_IN_B16),
		.SB_T1_NORTH_SB_OUT_B16(SB_ID0_3TRACKS_B16_PE_SB_T1_NORTH_SB_OUT_B16),
		.SB_T1_SOUTH_SB_IN_B16(SB_T1_SOUTH_SB_IN_B16),
		.SB_T1_SOUTH_SB_OUT_B16(SB_ID0_3TRACKS_B16_PE_SB_T1_SOUTH_SB_OUT_B16),
		.SB_T1_WEST_SB_IN_B16(SB_T1_WEST_SB_IN_B16),
		.SB_T1_WEST_SB_OUT_B16(SB_ID0_3TRACKS_B16_PE_SB_T1_WEST_SB_OUT_B16),
		.SB_T2_EAST_SB_IN_B16(SB_T2_EAST_SB_IN_B16),
		.SB_T2_EAST_SB_OUT_B16(SB_ID0_3TRACKS_B16_PE_SB_T2_EAST_SB_OUT_B16),
		.SB_T2_NORTH_SB_IN_B16(SB_T2_NORTH_SB_IN_B16),
		.SB_T2_NORTH_SB_OUT_B16(SB_ID0_3TRACKS_B16_PE_SB_T2_NORTH_SB_OUT_B16),
		.SB_T2_SOUTH_SB_IN_B16(SB_T2_SOUTH_SB_IN_B16),
		.SB_T2_SOUTH_SB_OUT_B16(SB_ID0_3TRACKS_B16_PE_SB_T2_SOUTH_SB_OUT_B16),
		.SB_T2_WEST_SB_IN_B16(SB_T2_WEST_SB_IN_B16),
		.SB_T2_WEST_SB_OUT_B16(SB_ID0_3TRACKS_B16_PE_SB_T2_WEST_SB_OUT_B16),
		.alu_res(PE_inst0_alu_res),
		.clk(clk),
		.config_config_addr(SB_ID0_3TRACKS_B16_PE_config_config_addr_in),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_7_out),
		.read_config_data(SB_ID0_3TRACKS_B16_PE_read_config_data),
		.reset(reset),
		.stall(stall)
	);
	mantle_wire__typeBitIn8 SB_ID0_3TRACKS_B16_PE_config_config_addr(
		.in(SB_ID0_3TRACKS_B16_PE_config_config_addr_in),
		.out(self_config_config_addr_out[31:24])
	);
	SB_ID0_3TRACKS_B1_PE SB_ID0_3TRACKS_B1_PE(
		.SB_T0_EAST_SB_IN_B1(SB_T0_EAST_SB_IN_B1),
		.SB_T0_EAST_SB_OUT_B1(SB_ID0_3TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_NORTH_SB_IN_B1(SB_T0_NORTH_SB_IN_B1),
		.SB_T0_NORTH_SB_OUT_B1(SB_ID0_3TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_IN_B1(SB_T0_SOUTH_SB_IN_B1),
		.SB_T0_SOUTH_SB_OUT_B1(SB_ID0_3TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_WEST_SB_IN_B1(SB_T0_WEST_SB_IN_B1),
		.SB_T0_WEST_SB_OUT_B1(SB_ID0_3TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1),
		.SB_T1_EAST_SB_IN_B1(SB_T1_EAST_SB_IN_B1),
		.SB_T1_EAST_SB_OUT_B1(SB_ID0_3TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_NORTH_SB_IN_B1(SB_T1_NORTH_SB_IN_B1),
		.SB_T1_NORTH_SB_OUT_B1(SB_ID0_3TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_IN_B1(SB_T1_SOUTH_SB_IN_B1),
		.SB_T1_SOUTH_SB_OUT_B1(SB_ID0_3TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_WEST_SB_IN_B1(SB_T1_WEST_SB_IN_B1),
		.SB_T1_WEST_SB_OUT_B1(SB_ID0_3TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1),
		.SB_T2_EAST_SB_IN_B1(SB_T2_EAST_SB_IN_B1),
		.SB_T2_EAST_SB_OUT_B1(SB_ID0_3TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_NORTH_SB_IN_B1(SB_T2_NORTH_SB_IN_B1),
		.SB_T2_NORTH_SB_OUT_B1(SB_ID0_3TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_IN_B1(SB_T2_SOUTH_SB_IN_B1),
		.SB_T2_SOUTH_SB_OUT_B1(SB_ID0_3TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_WEST_SB_IN_B1(SB_T2_WEST_SB_IN_B1),
		.SB_T2_WEST_SB_OUT_B1(SB_ID0_3TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1),
		.clk(clk),
		.config_config_addr(SB_ID0_3TRACKS_B1_PE_config_config_addr_in),
		.config_config_data(config_config_data),
		.config_read(config_read),
		.config_write(FEATURE_AND_6_out),
		.read_config_data(SB_ID0_3TRACKS_B1_PE_read_config_data),
		.res_p(PE_inst0_res_p),
		.reset(reset),
		.stall(stall)
	);
	mantle_wire__typeBitIn8 SB_ID0_3TRACKS_B1_PE_config_config_addr(
		.in(SB_ID0_3TRACKS_B1_PE_config_config_addr_in),
		.out(self_config_config_addr_out[31:24])
	);
	MuxWrapper_1_1 WIRE_SB_T0_EAST_SB_IN_B1(
		.I(SB_T0_EAST_SB_IN_B1),
		.O(WIRE_SB_T0_EAST_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T0_EAST_SB_IN_B16(
		.I(SB_T0_EAST_SB_IN_B16),
		.O(WIRE_SB_T0_EAST_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T0_NORTH_SB_IN_B1(
		.I(SB_T0_NORTH_SB_IN_B1),
		.O(WIRE_SB_T0_NORTH_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T0_NORTH_SB_IN_B16(
		.I(SB_T0_NORTH_SB_IN_B16),
		.O(WIRE_SB_T0_NORTH_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T0_SOUTH_SB_IN_B1(
		.I(SB_T0_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T0_SOUTH_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T0_SOUTH_SB_IN_B16(
		.I(SB_T0_SOUTH_SB_IN_B16),
		.O(WIRE_SB_T0_SOUTH_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T0_WEST_SB_IN_B1(
		.I(SB_T0_WEST_SB_IN_B1),
		.O(WIRE_SB_T0_WEST_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T0_WEST_SB_IN_B16(
		.I(SB_T0_WEST_SB_IN_B16),
		.O(WIRE_SB_T0_WEST_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T1_EAST_SB_IN_B1(
		.I(SB_T1_EAST_SB_IN_B1),
		.O(WIRE_SB_T1_EAST_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T1_EAST_SB_IN_B16(
		.I(SB_T1_EAST_SB_IN_B16),
		.O(WIRE_SB_T1_EAST_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T1_NORTH_SB_IN_B1(
		.I(SB_T1_NORTH_SB_IN_B1),
		.O(WIRE_SB_T1_NORTH_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T1_NORTH_SB_IN_B16(
		.I(SB_T1_NORTH_SB_IN_B16),
		.O(WIRE_SB_T1_NORTH_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T1_SOUTH_SB_IN_B1(
		.I(SB_T1_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T1_SOUTH_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T1_SOUTH_SB_IN_B16(
		.I(SB_T1_SOUTH_SB_IN_B16),
		.O(WIRE_SB_T1_SOUTH_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T1_WEST_SB_IN_B1(
		.I(SB_T1_WEST_SB_IN_B1),
		.O(WIRE_SB_T1_WEST_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T1_WEST_SB_IN_B16(
		.I(SB_T1_WEST_SB_IN_B16),
		.O(WIRE_SB_T1_WEST_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T2_EAST_SB_IN_B1(
		.I(SB_T2_EAST_SB_IN_B1),
		.O(WIRE_SB_T2_EAST_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T2_EAST_SB_IN_B16(
		.I(SB_T2_EAST_SB_IN_B16),
		.O(WIRE_SB_T2_EAST_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T2_NORTH_SB_IN_B1(
		.I(SB_T2_NORTH_SB_IN_B1),
		.O(WIRE_SB_T2_NORTH_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T2_NORTH_SB_IN_B16(
		.I(SB_T2_NORTH_SB_IN_B16),
		.O(WIRE_SB_T2_NORTH_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T2_SOUTH_SB_IN_B1(
		.I(SB_T2_SOUTH_SB_IN_B1),
		.O(WIRE_SB_T2_SOUTH_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T2_SOUTH_SB_IN_B16(
		.I(SB_T2_SOUTH_SB_IN_B16),
		.O(WIRE_SB_T2_SOUTH_SB_IN_B16_O)
	);
	MuxWrapper_1_1 WIRE_SB_T2_WEST_SB_IN_B1(
		.I(SB_T2_WEST_SB_IN_B1),
		.O(WIRE_SB_T2_WEST_SB_IN_B1_O)
	);
	MuxWrapper_1_16 WIRE_SB_T2_WEST_SB_IN_B16(
		.I(SB_T2_WEST_SB_IN_B16),
		.O(WIRE_SB_T2_WEST_SB_IN_B16_O)
	);
	corebit_and and_inst0(
		.in0(coreir_eq_16_inst0_out),
		.in1(config_read[0]),
		.out(and_inst0_out)
	);
	corebit_and and_inst1(
		.in0(coreir_eq_16_inst0_out),
		.in1(config_write[0]),
		.out(and_inst1_out)
	);
	coreir_const #(
		.value(8'h00),
		.width(8)
	) const_0_8(.out(const_0_8_out));
	coreir_const #(
		.value(9'h1ff),
		.width(9)
	) const_511_9(.out(const_511_9_out));
	coreir_eq #(.width(16)) coreir_eq_16_inst0(
		.in0(tile_id),
		.in1(self_config_config_addr_out[15:0]),
		.out(coreir_eq_16_inst0_out)
	);
	coreir_or #(.width(32)) read_config_data_or_inst0(
		.in0(read_data_mux_O),
		.in1(read_config_data_in),
		.out(read_config_data_or_inst0_out)
	);
	MuxWithDefaultWrapper_8_32_8_0 read_data_mux(
		.EN(and_inst0_out),
		.I_0(PE_inst0_read_config_data),
		.I_1(CB_bit0_read_config_data),
		.I_2(CB_bit1_read_config_data),
		.I_3(CB_bit2_read_config_data),
		.I_4(CB_data0_read_config_data),
		.I_5(CB_data1_read_config_data),
		.I_6(SB_ID0_3TRACKS_B1_PE_read_config_data),
		.I_7(SB_ID0_3TRACKS_B16_PE_read_config_data),
		.O(read_data_mux_O),
		.S(read_data_mux_S_in)
	);
	mantle_wire__typeBitIn8 read_data_mux_S(
		.in(read_data_mux_S_in),
		.out(self_config_config_addr_out[23:16])
	);
	mantle_wire__typeBit32 self_config_config_addr(
		.in(config_config_addr),
		.out(self_config_config_addr_out)
	);
	assign SB_T0_EAST_SB_OUT_B1 = SB_ID0_3TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1;
	assign SB_T0_EAST_SB_OUT_B16 = SB_ID0_3TRACKS_B16_PE_SB_T0_EAST_SB_OUT_B16;
	assign SB_T0_NORTH_SB_OUT_B1 = SB_ID0_3TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1;
	assign SB_T0_NORTH_SB_OUT_B16 = SB_ID0_3TRACKS_B16_PE_SB_T0_NORTH_SB_OUT_B16;
	assign SB_T0_SOUTH_SB_OUT_B1 = SB_ID0_3TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1;
	assign SB_T0_SOUTH_SB_OUT_B16 = SB_ID0_3TRACKS_B16_PE_SB_T0_SOUTH_SB_OUT_B16;
	assign SB_T0_WEST_SB_OUT_B1 = SB_ID0_3TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1;
	assign SB_T0_WEST_SB_OUT_B16 = SB_ID0_3TRACKS_B16_PE_SB_T0_WEST_SB_OUT_B16;
	assign SB_T1_EAST_SB_OUT_B1 = SB_ID0_3TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1;
	assign SB_T1_EAST_SB_OUT_B16 = SB_ID0_3TRACKS_B16_PE_SB_T1_EAST_SB_OUT_B16;
	assign SB_T1_NORTH_SB_OUT_B1 = SB_ID0_3TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1;
	assign SB_T1_NORTH_SB_OUT_B16 = SB_ID0_3TRACKS_B16_PE_SB_T1_NORTH_SB_OUT_B16;
	assign SB_T1_SOUTH_SB_OUT_B1 = SB_ID0_3TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1;
	assign SB_T1_SOUTH_SB_OUT_B16 = SB_ID0_3TRACKS_B16_PE_SB_T1_SOUTH_SB_OUT_B16;
	assign SB_T1_WEST_SB_OUT_B1 = SB_ID0_3TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1;
	assign SB_T1_WEST_SB_OUT_B16 = SB_ID0_3TRACKS_B16_PE_SB_T1_WEST_SB_OUT_B16;
	assign SB_T2_EAST_SB_OUT_B1 = SB_ID0_3TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1;
	assign SB_T2_EAST_SB_OUT_B16 = SB_ID0_3TRACKS_B16_PE_SB_T2_EAST_SB_OUT_B16;
	assign SB_T2_NORTH_SB_OUT_B1 = SB_ID0_3TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1;
	assign SB_T2_NORTH_SB_OUT_B16 = SB_ID0_3TRACKS_B16_PE_SB_T2_NORTH_SB_OUT_B16;
	assign SB_T2_SOUTH_SB_OUT_B1 = SB_ID0_3TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1;
	assign SB_T2_SOUTH_SB_OUT_B16 = SB_ID0_3TRACKS_B16_PE_SB_T2_SOUTH_SB_OUT_B16;
	assign SB_T2_WEST_SB_OUT_B1 = SB_ID0_3TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1;
	assign SB_T2_WEST_SB_OUT_B16 = SB_ID0_3TRACKS_B16_PE_SB_T2_WEST_SB_OUT_B16;
	assign clk_out = clk_pass_through;
	assign clk_pass_through_out_bot = clk_pass_through;
	assign config_out_config_addr = config_config_addr;
	assign config_out_config_data = config_config_data;
	assign config_out_read = config_read;
	assign config_out_write = config_write;
	assign hi = const_511_9_out;
	assign lo = const_0_8_out;
	assign read_config_data = read_config_data_or_inst0_out;
	assign reset_out = reset;
	assign stall_out = stall;
endmodule
module Interconnect (
	clk,
	config_0_config_addr,
	config_0_config_data,
	config_0_read,
	config_0_write,
	config_1_config_addr,
	config_1_config_data,
	config_1_read,
	config_1_write,
	config_2_config_addr,
	config_2_config_data,
	config_2_read,
	config_2_write,
	config_3_config_addr,
	config_3_config_data,
	config_3_read,
	config_3_write,
	glb2io_16_X00_Y00,
	glb2io_16_X01_Y00,
	// glb2io_16_X02_Y00,
	// glb2io_16_X03_Y00,
	glb2io_1_X00_Y00,
	glb2io_1_X01_Y00,
	// glb2io_1_X02_Y00,
	// glb2io_1_X03_Y00,
	io2glb_16_X00_Y00,
	io2glb_16_X01_Y00,
	// io2glb_16_X02_Y00,
	// io2glb_16_X03_Y00,
	io2glb_1_X00_Y00,
	io2glb_1_X01_Y00,
	// io2glb_1_X02_Y00,
	// io2glb_1_X03_Y00,
	read_config_data,
	reset,
	stall
);
	input clk;
	input [31:0] config_0_config_addr;
	input [31:0] config_0_config_data;
	input [0:0] config_0_read;
	input [0:0] config_0_write;
	input [31:0] config_1_config_addr;
	input [31:0] config_1_config_data;
	input [0:0] config_1_read;
	input [0:0] config_1_write;
	input [31:0] config_2_config_addr;
	input [31:0] config_2_config_data;
	input [0:0] config_2_read;
	input [0:0] config_2_write;
	input [31:0] config_3_config_addr;
	input [31:0] config_3_config_data;
	input [0:0] config_3_read;
	input [0:0] config_3_write;
	input [15:0] glb2io_16_X00_Y00;
	input [15:0] glb2io_16_X01_Y00;
	// input [15:0] glb2io_16_X02_Y00;
	// input [15:0] glb2io_16_X03_Y00;
	input [0:0] glb2io_1_X00_Y00;
	input [0:0] glb2io_1_X01_Y00;
	// input [0:0] glb2io_1_X02_Y00;
	// input [0:0] glb2io_1_X03_Y00;
	output [15:0] io2glb_16_X00_Y00;
	output [15:0] io2glb_16_X01_Y00;
	// output [15:0] io2glb_16_X02_Y00;
	// output [15:0] io2glb_16_X03_Y00;
	output [0:0] io2glb_1_X00_Y00;
	output [0:0] io2glb_1_X01_Y00;
	// output [0:0] io2glb_1_X02_Y00;
	// output [0:0] io2glb_1_X03_Y00;
	output [31:0] read_config_data;
	input reset;
	input [3:0] stall;
	wire [0:0] Tile_X00_Y00_io2glb_1;
	wire [0:0] Tile_X00_Y00_io2f_1;
	wire [15:0] Tile_X00_Y00_io2glb_16;
	wire [15:0] Tile_X00_Y00_io2f_16;
	wire [8:0] Tile_X00_Y00_hi;
	wire [7:0] Tile_X00_Y00_lo;
	wire [0:0] Tile_X00_Y01_SB_T0_EAST_SB_OUT_B1;
	wire [15:0] Tile_X00_Y01_SB_T0_EAST_SB_OUT_B16;
	wire [0:0] Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B1;
	wire [15:0] Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B16;
	wire [0:0] Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B1;
	wire [15:0] Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B16;
	wire [0:0] Tile_X00_Y01_SB_T0_WEST_SB_OUT_B1;
	wire [15:0] Tile_X00_Y01_SB_T0_WEST_SB_OUT_B16;
	wire [0:0] Tile_X00_Y01_SB_T1_EAST_SB_OUT_B1;
	wire [15:0] Tile_X00_Y01_SB_T1_EAST_SB_OUT_B16;
	wire [0:0] Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B1;
	wire [15:0] Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B16;
	wire [0:0] Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B1;
	wire [15:0] Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B16;
	wire [0:0] Tile_X00_Y01_SB_T1_WEST_SB_OUT_B1;
	wire [15:0] Tile_X00_Y01_SB_T1_WEST_SB_OUT_B16;
	wire [0:0] Tile_X00_Y01_SB_T2_EAST_SB_OUT_B1;
	wire [15:0] Tile_X00_Y01_SB_T2_EAST_SB_OUT_B16;
	wire [0:0] Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B1;
	wire [15:0] Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B16;
	wire [0:0] Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B1;
	wire [15:0] Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B16;
	wire [0:0] Tile_X00_Y01_SB_T2_WEST_SB_OUT_B1;
	wire [15:0] Tile_X00_Y01_SB_T2_WEST_SB_OUT_B16;
	wire Tile_X00_Y01_clk_out;
	wire Tile_X00_Y01_clk_pass_through_out_bot;
	wire [31:0] Tile_X00_Y01_config_out_config_addr;
	wire [31:0] Tile_X00_Y01_config_out_config_data;
	wire [0:0] Tile_X00_Y01_config_out_read;
	wire [0:0] Tile_X00_Y01_config_out_write;
	wire [8:0] Tile_X00_Y01_hi;
	wire [7:0] Tile_X00_Y01_lo_unq1;
	wire [31:0] Tile_X00_Y01_read_config_data;
	wire Tile_X00_Y01_reset_out;
	wire [0:0] Tile_X00_Y01_stall_out;
	wire [7:0] Tile_X00_Y01_lo_out;
	wire [15:0] Tile_X00_Y01_tile_id_in;
	wire [0:0] Tile_X00_Y02_SB_T0_EAST_SB_OUT_B1;
	wire [15:0] Tile_X00_Y02_SB_T0_EAST_SB_OUT_B16;
	wire [0:0] Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B1;
	wire [15:0] Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B16;
	wire [0:0] Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B1;
	wire [15:0] Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B16;
	wire [0:0] Tile_X00_Y02_SB_T0_WEST_SB_OUT_B1;
	wire [15:0] Tile_X00_Y02_SB_T0_WEST_SB_OUT_B16;
	wire [0:0] Tile_X00_Y02_SB_T1_EAST_SB_OUT_B1;
	wire [15:0] Tile_X00_Y02_SB_T1_EAST_SB_OUT_B16;
	wire [0:0] Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B1;
	wire [15:0] Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B16;
	wire [0:0] Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B1;
	wire [15:0] Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B16;
	wire [0:0] Tile_X00_Y02_SB_T1_WEST_SB_OUT_B1;
	wire [15:0] Tile_X00_Y02_SB_T1_WEST_SB_OUT_B16;
	wire [0:0] Tile_X00_Y02_SB_T2_EAST_SB_OUT_B1;
	wire [15:0] Tile_X00_Y02_SB_T2_EAST_SB_OUT_B16;
	wire [0:0] Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B1;
	wire [15:0] Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B16;
	wire [0:0] Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B1;
	wire [15:0] Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B16;
	wire [0:0] Tile_X00_Y02_SB_T2_WEST_SB_OUT_B1;
	wire [15:0] Tile_X00_Y02_SB_T2_WEST_SB_OUT_B16;
	wire Tile_X00_Y02_clk_out;
	wire Tile_X00_Y02_clk_pass_through_out_bot;
	wire [31:0] Tile_X00_Y02_config_out_config_addr;
	wire [31:0] Tile_X00_Y02_config_out_config_data;
	wire [0:0] Tile_X00_Y02_config_out_read;
	wire [0:0] Tile_X00_Y02_config_out_write;
	wire [8:0] Tile_X00_Y02_hi;
	wire [7:0] Tile_X00_Y02_lo_unq1;
	wire [31:0] Tile_X00_Y02_read_config_data;
	wire Tile_X00_Y02_reset_out;
	wire [0:0] Tile_X00_Y02_stall_out;
	wire [7:0] Tile_X00_Y02_lo_out;
	wire [15:0] Tile_X00_Y02_tile_id_in;
	// wire [0:0] Tile_X00_Y03_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y03_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y03_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y03_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y03_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y03_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y03_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y03_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y03_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y03_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y03_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y03_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X00_Y03_clk_out;
	// wire Tile_X00_Y03_clk_pass_through_out_bot;
	// wire [31:0] Tile_X00_Y03_config_out_config_addr;
	// wire [31:0] Tile_X00_Y03_config_out_config_data;
	// wire [0:0] Tile_X00_Y03_config_out_read;
	// wire [0:0] Tile_X00_Y03_config_out_write;
	// wire [8:0] Tile_X00_Y03_hi_unq1;
	// wire [7:0] Tile_X00_Y03_lo_unq1;
	// wire [31:0] Tile_X00_Y03_read_config_data;
	// wire Tile_X00_Y03_reset_out;
	// wire [0:0] Tile_X00_Y03_stall_out;
	// wire [8:0] Tile_X00_Y03_hi_out;
	// wire [7:0] Tile_X00_Y03_lo_out;
	// wire [15:0] Tile_X00_Y03_tile_id_in;
	// wire [0:0] Tile_X00_Y04_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y04_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y04_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y04_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y04_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y04_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y04_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y04_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y04_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y04_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y04_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y04_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X00_Y04_clk_out;
	// wire Tile_X00_Y04_clk_pass_through_out_bot;
	// wire [31:0] Tile_X00_Y04_config_out_config_addr;
	// wire [31:0] Tile_X00_Y04_config_out_config_data;
	// wire [0:0] Tile_X00_Y04_config_out_read;
	// wire [0:0] Tile_X00_Y04_config_out_write;
	// wire [8:0] Tile_X00_Y04_hi;
	// wire [7:0] Tile_X00_Y04_lo_unq1;
	// wire [31:0] Tile_X00_Y04_read_config_data;
	// wire Tile_X00_Y04_reset_out;
	// wire [0:0] Tile_X00_Y04_stall_out;
	// wire [7:0] Tile_X00_Y04_lo_out;
	// wire [15:0] Tile_X00_Y04_tile_id_in;
	// wire [0:0] Tile_X00_Y05_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y05_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y05_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y05_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y05_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y05_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y05_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y05_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y05_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y05_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y05_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y05_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y05_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y05_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y05_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y05_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y05_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y05_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y05_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y05_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y05_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y05_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y05_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y05_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X00_Y05_clk_out;
	// wire Tile_X00_Y05_clk_pass_through_out_bot;
	// wire [31:0] Tile_X00_Y05_config_out_config_addr;
	// wire [31:0] Tile_X00_Y05_config_out_config_data;
	// wire [0:0] Tile_X00_Y05_config_out_read;
	// wire [0:0] Tile_X00_Y05_config_out_write;
	// wire [8:0] Tile_X00_Y05_hi;
	// wire [7:0] Tile_X00_Y05_lo_unq1;
	// wire [31:0] Tile_X00_Y05_read_config_data;
	// wire Tile_X00_Y05_reset_out;
	// wire [0:0] Tile_X00_Y05_stall_out;
	// wire [7:0] Tile_X00_Y05_lo_out;
	// wire [15:0] Tile_X00_Y05_tile_id_in;
	// wire [0:0] Tile_X00_Y06_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y06_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y06_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y06_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y06_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y06_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y06_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y06_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y06_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y06_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y06_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y06_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y06_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y06_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y06_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y06_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y06_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y06_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y06_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y06_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y06_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y06_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y06_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y06_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X00_Y06_clk_out;
	// wire Tile_X00_Y06_clk_pass_through_out_bot;
	// wire [31:0] Tile_X00_Y06_config_out_config_addr;
	// wire [31:0] Tile_X00_Y06_config_out_config_data;
	// wire [0:0] Tile_X00_Y06_config_out_read;
	// wire [0:0] Tile_X00_Y06_config_out_write;
	// wire [8:0] Tile_X00_Y06_hi;
	// wire [7:0] Tile_X00_Y06_lo_unq1;
	// wire [31:0] Tile_X00_Y06_read_config_data;
	// wire Tile_X00_Y06_reset_out;
	// wire [0:0] Tile_X00_Y06_stall_out;
	// wire [7:0] Tile_X00_Y06_lo_out;
	// wire [15:0] Tile_X00_Y06_tile_id_in;
	// wire [0:0] Tile_X00_Y07_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y07_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y07_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y07_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y07_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y07_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y07_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y07_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y07_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y07_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y07_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y07_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y07_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y07_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y07_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y07_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y07_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y07_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y07_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y07_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y07_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y07_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y07_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y07_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X00_Y07_clk_out;
	// wire Tile_X00_Y07_clk_pass_through_out_bot;
	// wire [31:0] Tile_X00_Y07_config_out_config_addr;
	// wire [31:0] Tile_X00_Y07_config_out_config_data;
	// wire [0:0] Tile_X00_Y07_config_out_read;
	// wire [0:0] Tile_X00_Y07_config_out_write;
	// wire [8:0] Tile_X00_Y07_hi_unq1;
	// wire [7:0] Tile_X00_Y07_lo_unq1;
	// wire [31:0] Tile_X00_Y07_read_config_data;
	// wire Tile_X00_Y07_reset_out;
	// wire [0:0] Tile_X00_Y07_stall_out;
	// wire [8:0] Tile_X00_Y07_hi_out;
	// wire [7:0] Tile_X00_Y07_lo_out;
	// wire [15:0] Tile_X00_Y07_tile_id_in;
	// wire [0:0] Tile_X00_Y08_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y08_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y08_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y08_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y08_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y08_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y08_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y08_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y08_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y08_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y08_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y08_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y08_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y08_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y08_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y08_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y08_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y08_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y08_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y08_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y08_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y08_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X00_Y08_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X00_Y08_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X00_Y08_clk_out;
	// wire Tile_X00_Y08_clk_pass_through_out_bot;
	// wire [31:0] Tile_X00_Y08_config_out_config_addr;
	// wire [31:0] Tile_X00_Y08_config_out_config_data;
	// wire [0:0] Tile_X00_Y08_config_out_read;
	// wire [0:0] Tile_X00_Y08_config_out_write;
	// wire [8:0] Tile_X00_Y08_hi;
	// wire [7:0] Tile_X00_Y08_lo_unq1;
	// wire [31:0] Tile_X00_Y08_read_config_data;
	// wire Tile_X00_Y08_reset_out;
	// wire [0:0] Tile_X00_Y08_stall_out;
	// wire [7:0] Tile_X00_Y08_lo_out;
	// wire [15:0] Tile_X00_Y08_tile_id_in;
	wire [0:0] Tile_X01_Y00_io2glb_1;
	wire [0:0] Tile_X01_Y00_io2f_1;
	wire [15:0] Tile_X01_Y00_io2glb_16;
	wire [15:0] Tile_X01_Y00_io2f_16;
	wire [8:0] Tile_X01_Y00_hi;
	wire [7:0] Tile_X01_Y00_lo;
	wire [0:0] Tile_X01_Y01_SB_T0_EAST_SB_OUT_B1;
	wire [15:0] Tile_X01_Y01_SB_T0_EAST_SB_OUT_B16;
	wire [0:0] Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B1;
	wire [15:0] Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B16;
	wire [0:0] Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B1;
	wire [15:0] Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B16;
	wire [0:0] Tile_X01_Y01_SB_T0_WEST_SB_OUT_B1;
	wire [15:0] Tile_X01_Y01_SB_T0_WEST_SB_OUT_B16;
	wire [0:0] Tile_X01_Y01_SB_T1_EAST_SB_OUT_B1;
	wire [15:0] Tile_X01_Y01_SB_T1_EAST_SB_OUT_B16;
	wire [0:0] Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B1;
	wire [15:0] Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B16;
	wire [0:0] Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B1;
	wire [15:0] Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B16;
	wire [0:0] Tile_X01_Y01_SB_T1_WEST_SB_OUT_B1;
	wire [15:0] Tile_X01_Y01_SB_T1_WEST_SB_OUT_B16;
	wire [0:0] Tile_X01_Y01_SB_T2_EAST_SB_OUT_B1;
	wire [15:0] Tile_X01_Y01_SB_T2_EAST_SB_OUT_B16;
	wire [0:0] Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B1;
	wire [15:0] Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B16;
	wire [0:0] Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B1;
	wire [15:0] Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B16;
	wire [0:0] Tile_X01_Y01_SB_T2_WEST_SB_OUT_B1;
	wire [15:0] Tile_X01_Y01_SB_T2_WEST_SB_OUT_B16;
	wire Tile_X01_Y01_clk_out;
	wire Tile_X01_Y01_clk_pass_through_out_bot;
	wire [31:0] Tile_X01_Y01_config_out_config_addr;
	wire [31:0] Tile_X01_Y01_config_out_config_data;
	wire [0:0] Tile_X01_Y01_config_out_read;
	wire [0:0] Tile_X01_Y01_config_out_write;
	wire [8:0] Tile_X01_Y01_hi;
	wire [7:0] Tile_X01_Y01_lo_unq1;
	wire [31:0] Tile_X01_Y01_read_config_data;
	wire Tile_X01_Y01_reset_out;
	wire [0:0] Tile_X01_Y01_stall_out;
	wire [7:0] Tile_X01_Y01_lo_out;
	wire [15:0] Tile_X01_Y01_tile_id_in;
	wire [0:0] Tile_X01_Y02_SB_T0_EAST_SB_OUT_B1;
	wire [15:0] Tile_X01_Y02_SB_T0_EAST_SB_OUT_B16;
	wire [0:0] Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B1;
	wire [15:0] Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B16;
	wire [0:0] Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B1;
	wire [15:0] Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B16;
	wire [0:0] Tile_X01_Y02_SB_T0_WEST_SB_OUT_B1;
	wire [15:0] Tile_X01_Y02_SB_T0_WEST_SB_OUT_B16;
	wire [0:0] Tile_X01_Y02_SB_T1_EAST_SB_OUT_B1;
	wire [15:0] Tile_X01_Y02_SB_T1_EAST_SB_OUT_B16;
	wire [0:0] Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B1;
	wire [15:0] Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B16;
	wire [0:0] Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B1;
	wire [15:0] Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B16;
	wire [0:0] Tile_X01_Y02_SB_T1_WEST_SB_OUT_B1;
	wire [15:0] Tile_X01_Y02_SB_T1_WEST_SB_OUT_B16;
	wire [0:0] Tile_X01_Y02_SB_T2_EAST_SB_OUT_B1;
	wire [15:0] Tile_X01_Y02_SB_T2_EAST_SB_OUT_B16;
	wire [0:0] Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B1;
	wire [15:0] Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B16;
	wire [0:0] Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B1;
	wire [15:0] Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B16;
	wire [0:0] Tile_X01_Y02_SB_T2_WEST_SB_OUT_B1;
	wire [15:0] Tile_X01_Y02_SB_T2_WEST_SB_OUT_B16;
	wire Tile_X01_Y02_clk_out;
	wire Tile_X01_Y02_clk_pass_through_out_bot;
	wire [31:0] Tile_X01_Y02_config_out_config_addr;
	wire [31:0] Tile_X01_Y02_config_out_config_data;
	wire [0:0] Tile_X01_Y02_config_out_read;
	wire [0:0] Tile_X01_Y02_config_out_write;
	wire [8:0] Tile_X01_Y02_hi;
	wire [7:0] Tile_X01_Y02_lo_unq1;
	wire [31:0] Tile_X01_Y02_read_config_data;
	wire Tile_X01_Y02_reset_out;
	wire [0:0] Tile_X01_Y02_stall_out;
	wire [7:0] Tile_X01_Y02_lo_out;
	wire [15:0] Tile_X01_Y02_tile_id_in;
	// wire [0:0] Tile_X01_Y03_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y03_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y03_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y03_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y03_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y03_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y03_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y03_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y03_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y03_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y03_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y03_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X01_Y03_clk_out;
	// wire Tile_X01_Y03_clk_pass_through_out_bot;
	// wire [31:0] Tile_X01_Y03_config_out_config_addr;
	// wire [31:0] Tile_X01_Y03_config_out_config_data;
	// wire [0:0] Tile_X01_Y03_config_out_read;
	// wire [0:0] Tile_X01_Y03_config_out_write;
	// wire [8:0] Tile_X01_Y03_hi_unq1;
	// wire [7:0] Tile_X01_Y03_lo_unq1;
	// wire [31:0] Tile_X01_Y03_read_config_data;
	// wire Tile_X01_Y03_reset_out;
	// wire [0:0] Tile_X01_Y03_stall_out;
	// wire [8:0] Tile_X01_Y03_hi_out;
	// wire [7:0] Tile_X01_Y03_lo_out;
	// wire [15:0] Tile_X01_Y03_tile_id_in;
	// wire [0:0] Tile_X01_Y04_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y04_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y04_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y04_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y04_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y04_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y04_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y04_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y04_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y04_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y04_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y04_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X01_Y04_clk_out;
	// wire Tile_X01_Y04_clk_pass_through_out_bot;
	// wire [31:0] Tile_X01_Y04_config_out_config_addr;
	// wire [31:0] Tile_X01_Y04_config_out_config_data;
	// wire [0:0] Tile_X01_Y04_config_out_read;
	// wire [0:0] Tile_X01_Y04_config_out_write;
	// wire [8:0] Tile_X01_Y04_hi;
	// wire [7:0] Tile_X01_Y04_lo_unq1;
	// wire [31:0] Tile_X01_Y04_read_config_data;
	// wire Tile_X01_Y04_reset_out;
	// wire [0:0] Tile_X01_Y04_stall_out;
	// wire [7:0] Tile_X01_Y04_lo_out;
	// wire [15:0] Tile_X01_Y04_tile_id_in;
	// wire [0:0] Tile_X01_Y05_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y05_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y05_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y05_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y05_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y05_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y05_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y05_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y05_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y05_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y05_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y05_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y05_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y05_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y05_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y05_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y05_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y05_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y05_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y05_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y05_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y05_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y05_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y05_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X01_Y05_clk_out;
	// wire Tile_X01_Y05_clk_pass_through_out_bot;
	// wire [31:0] Tile_X01_Y05_config_out_config_addr;
	// wire [31:0] Tile_X01_Y05_config_out_config_data;
	// wire [0:0] Tile_X01_Y05_config_out_read;
	// wire [0:0] Tile_X01_Y05_config_out_write;
	// wire [8:0] Tile_X01_Y05_hi;
	// wire [7:0] Tile_X01_Y05_lo_unq1;
	// wire [31:0] Tile_X01_Y05_read_config_data;
	// wire Tile_X01_Y05_reset_out;
	// wire [0:0] Tile_X01_Y05_stall_out;
	// wire [7:0] Tile_X01_Y05_lo_out;
	// wire [15:0] Tile_X01_Y05_tile_id_in;
	// wire [0:0] Tile_X01_Y06_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y06_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y06_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y06_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y06_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y06_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y06_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y06_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y06_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y06_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y06_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y06_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y06_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y06_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y06_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y06_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y06_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y06_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y06_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y06_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y06_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y06_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y06_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y06_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X01_Y06_clk_out;
	// wire Tile_X01_Y06_clk_pass_through_out_bot;
	// wire [31:0] Tile_X01_Y06_config_out_config_addr;
	// wire [31:0] Tile_X01_Y06_config_out_config_data;
	// wire [0:0] Tile_X01_Y06_config_out_read;
	// wire [0:0] Tile_X01_Y06_config_out_write;
	// wire [8:0] Tile_X01_Y06_hi;
	// wire [7:0] Tile_X01_Y06_lo_unq1;
	// wire [31:0] Tile_X01_Y06_read_config_data;
	// wire Tile_X01_Y06_reset_out;
	// wire [0:0] Tile_X01_Y06_stall_out;
	// wire [7:0] Tile_X01_Y06_lo_out;
	// wire [15:0] Tile_X01_Y06_tile_id_in;
	// wire [0:0] Tile_X01_Y07_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y07_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y07_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y07_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y07_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y07_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y07_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y07_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y07_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y07_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y07_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y07_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y07_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y07_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y07_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y07_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y07_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y07_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y07_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y07_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y07_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y07_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y07_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y07_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X01_Y07_clk_out;
	// wire Tile_X01_Y07_clk_pass_through_out_bot;
	// wire [31:0] Tile_X01_Y07_config_out_config_addr;
	// wire [31:0] Tile_X01_Y07_config_out_config_data;
	// wire [0:0] Tile_X01_Y07_config_out_read;
	// wire [0:0] Tile_X01_Y07_config_out_write;
	// wire [8:0] Tile_X01_Y07_hi_unq1;
	// wire [7:0] Tile_X01_Y07_lo_unq1;
	// wire [31:0] Tile_X01_Y07_read_config_data;
	// wire Tile_X01_Y07_reset_out;
	// wire [0:0] Tile_X01_Y07_stall_out;
	// wire [8:0] Tile_X01_Y07_hi_out;
	// wire [7:0] Tile_X01_Y07_lo_out;
	// wire [15:0] Tile_X01_Y07_tile_id_in;
	// wire [0:0] Tile_X01_Y08_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y08_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y08_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y08_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y08_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y08_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y08_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y08_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y08_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y08_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y08_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y08_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y08_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y08_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y08_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y08_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y08_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y08_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y08_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y08_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y08_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y08_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X01_Y08_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X01_Y08_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X01_Y08_clk_out;
	// wire Tile_X01_Y08_clk_pass_through_out_bot;
	// wire [31:0] Tile_X01_Y08_config_out_config_addr;
	// wire [31:0] Tile_X01_Y08_config_out_config_data;
	// wire [0:0] Tile_X01_Y08_config_out_read;
	// wire [0:0] Tile_X01_Y08_config_out_write;
	// wire [8:0] Tile_X01_Y08_hi;
	// wire [7:0] Tile_X01_Y08_lo_unq1;
	// wire [31:0] Tile_X01_Y08_read_config_data;
	// wire Tile_X01_Y08_reset_out;
	// wire [0:0] Tile_X01_Y08_stall_out;
	// wire [7:0] Tile_X01_Y08_lo_out;
	// wire [15:0] Tile_X01_Y08_tile_id_in;
	// wire [0:0] Tile_X02_Y00_io2glb_1;
	// wire [0:0] Tile_X02_Y00_io2f_1;
	// wire [15:0] Tile_X02_Y00_io2glb_16;
	// wire [15:0] Tile_X02_Y00_io2f_16;
	// wire [8:0] Tile_X02_Y00_hi;
	// wire [7:0] Tile_X02_Y00_lo;
	// wire [0:0] Tile_X02_Y01_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y01_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y01_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y01_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y01_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y01_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y01_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y01_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y01_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y01_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y01_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y01_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X02_Y01_clk_out;
	// wire Tile_X02_Y01_clk_pass_through_out_bot;
	// wire [31:0] Tile_X02_Y01_config_out_config_addr;
	// wire [31:0] Tile_X02_Y01_config_out_config_data;
	// wire [0:0] Tile_X02_Y01_config_out_read;
	// wire [0:0] Tile_X02_Y01_config_out_write;
	// wire [8:0] Tile_X02_Y01_hi;
	// wire [7:0] Tile_X02_Y01_lo_unq1;
	// wire [31:0] Tile_X02_Y01_read_config_data;
	// wire Tile_X02_Y01_reset_out;
	// wire [0:0] Tile_X02_Y01_stall_out;
	// wire [7:0] Tile_X02_Y01_lo_out;
	// wire [15:0] Tile_X02_Y01_tile_id_in;
	// wire [0:0] Tile_X02_Y02_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y02_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y02_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y02_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y02_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y02_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y02_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y02_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y02_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y02_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y02_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y02_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X02_Y02_clk_out;
	// wire Tile_X02_Y02_clk_pass_through_out_bot;
	// wire [31:0] Tile_X02_Y02_config_out_config_addr;
	// wire [31:0] Tile_X02_Y02_config_out_config_data;
	// wire [0:0] Tile_X02_Y02_config_out_read;
	// wire [0:0] Tile_X02_Y02_config_out_write;
	// wire [8:0] Tile_X02_Y02_hi;
	// wire [7:0] Tile_X02_Y02_lo_unq1;
	// wire [31:0] Tile_X02_Y02_read_config_data;
	// wire Tile_X02_Y02_reset_out;
	// wire [0:0] Tile_X02_Y02_stall_out;
	// wire [7:0] Tile_X02_Y02_lo_out;
	// wire [15:0] Tile_X02_Y02_tile_id_in;
	// wire [0:0] Tile_X02_Y03_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y03_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y03_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y03_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y03_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y03_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y03_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y03_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y03_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y03_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y03_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y03_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X02_Y03_clk_out;
	// wire Tile_X02_Y03_clk_pass_through_out_bot;
	// wire [31:0] Tile_X02_Y03_config_out_config_addr;
	// wire [31:0] Tile_X02_Y03_config_out_config_data;
	// wire [0:0] Tile_X02_Y03_config_out_read;
	// wire [0:0] Tile_X02_Y03_config_out_write;
	// wire [8:0] Tile_X02_Y03_hi_unq1;
	// wire [7:0] Tile_X02_Y03_lo_unq1;
	// wire [31:0] Tile_X02_Y03_read_config_data;
	// wire Tile_X02_Y03_reset_out;
	// wire [0:0] Tile_X02_Y03_stall_out;
	// wire [8:0] Tile_X02_Y03_hi_out;
	// wire [7:0] Tile_X02_Y03_lo_out;
	// wire [15:0] Tile_X02_Y03_tile_id_in;
	// wire [0:0] Tile_X02_Y04_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y04_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y04_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y04_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y04_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y04_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y04_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y04_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y04_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y04_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y04_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y04_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X02_Y04_clk_out;
	// wire Tile_X02_Y04_clk_pass_through_out_bot;
	// wire [31:0] Tile_X02_Y04_config_out_config_addr;
	// wire [31:0] Tile_X02_Y04_config_out_config_data;
	// wire [0:0] Tile_X02_Y04_config_out_read;
	// wire [0:0] Tile_X02_Y04_config_out_write;
	// wire [8:0] Tile_X02_Y04_hi;
	// wire [7:0] Tile_X02_Y04_lo_unq1;
	// wire [31:0] Tile_X02_Y04_read_config_data;
	// wire Tile_X02_Y04_reset_out;
	// wire [0:0] Tile_X02_Y04_stall_out;
	// wire [7:0] Tile_X02_Y04_lo_out;
	// wire [15:0] Tile_X02_Y04_tile_id_in;
	// wire [0:0] Tile_X02_Y05_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y05_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y05_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y05_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y05_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y05_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y05_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y05_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y05_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y05_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y05_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y05_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y05_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y05_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y05_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y05_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y05_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y05_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y05_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y05_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y05_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y05_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y05_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y05_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X02_Y05_clk_out;
	// wire Tile_X02_Y05_clk_pass_through_out_bot;
	// wire [31:0] Tile_X02_Y05_config_out_config_addr;
	// wire [31:0] Tile_X02_Y05_config_out_config_data;
	// wire [0:0] Tile_X02_Y05_config_out_read;
	// wire [0:0] Tile_X02_Y05_config_out_write;
	// wire [8:0] Tile_X02_Y05_hi;
	// wire [7:0] Tile_X02_Y05_lo_unq1;
	// wire [31:0] Tile_X02_Y05_read_config_data;
	// wire Tile_X02_Y05_reset_out;
	// wire [0:0] Tile_X02_Y05_stall_out;
	// wire [7:0] Tile_X02_Y05_lo_out;
	// wire [15:0] Tile_X02_Y05_tile_id_in;
	// wire [0:0] Tile_X02_Y06_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y06_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y06_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y06_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y06_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y06_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y06_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y06_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y06_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y06_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y06_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y06_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y06_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y06_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y06_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y06_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y06_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y06_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y06_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y06_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y06_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y06_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y06_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y06_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X02_Y06_clk_out;
	// wire Tile_X02_Y06_clk_pass_through_out_bot;
	// wire [31:0] Tile_X02_Y06_config_out_config_addr;
	// wire [31:0] Tile_X02_Y06_config_out_config_data;
	// wire [0:0] Tile_X02_Y06_config_out_read;
	// wire [0:0] Tile_X02_Y06_config_out_write;
	// wire [8:0] Tile_X02_Y06_hi;
	// wire [7:0] Tile_X02_Y06_lo_unq1;
	// wire [31:0] Tile_X02_Y06_read_config_data;
	// wire Tile_X02_Y06_reset_out;
	// wire [0:0] Tile_X02_Y06_stall_out;
	// wire [7:0] Tile_X02_Y06_lo_out;
	// wire [15:0] Tile_X02_Y06_tile_id_in;
	// wire [0:0] Tile_X02_Y07_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y07_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y07_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y07_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y07_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y07_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y07_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y07_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y07_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y07_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y07_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y07_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y07_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y07_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y07_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y07_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y07_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y07_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y07_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y07_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y07_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y07_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y07_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y07_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X02_Y07_clk_out;
	// wire Tile_X02_Y07_clk_pass_through_out_bot;
	// wire [31:0] Tile_X02_Y07_config_out_config_addr;
	// wire [31:0] Tile_X02_Y07_config_out_config_data;
	// wire [0:0] Tile_X02_Y07_config_out_read;
	// wire [0:0] Tile_X02_Y07_config_out_write;
	// wire [8:0] Tile_X02_Y07_hi_unq1;
	// wire [7:0] Tile_X02_Y07_lo_unq1;
	// wire [31:0] Tile_X02_Y07_read_config_data;
	// wire Tile_X02_Y07_reset_out;
	// wire [0:0] Tile_X02_Y07_stall_out;
	// wire [8:0] Tile_X02_Y07_hi_out;
	// wire [7:0] Tile_X02_Y07_lo_out;
	// wire [15:0] Tile_X02_Y07_tile_id_in;
	// wire [0:0] Tile_X02_Y08_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y08_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y08_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y08_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y08_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y08_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y08_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y08_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y08_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y08_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y08_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y08_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y08_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y08_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y08_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y08_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y08_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y08_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y08_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y08_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y08_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y08_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X02_Y08_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X02_Y08_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X02_Y08_clk_out;
	// wire Tile_X02_Y08_clk_pass_through_out_bot;
	// wire [31:0] Tile_X02_Y08_config_out_config_addr;
	// wire [31:0] Tile_X02_Y08_config_out_config_data;
	// wire [0:0] Tile_X02_Y08_config_out_read;
	// wire [0:0] Tile_X02_Y08_config_out_write;
	// wire [8:0] Tile_X02_Y08_hi;
	// wire [7:0] Tile_X02_Y08_lo_unq1;
	// wire [31:0] Tile_X02_Y08_read_config_data;
	// wire Tile_X02_Y08_reset_out;
	// wire [0:0] Tile_X02_Y08_stall_out;
	// wire [7:0] Tile_X02_Y08_lo_out;
	// wire [15:0] Tile_X02_Y08_tile_id_in;
	// wire [0:0] Tile_X03_Y00_io2glb_1;
	// wire [0:0] Tile_X03_Y00_io2f_1;
	// wire [15:0] Tile_X03_Y00_io2glb_16;
	// wire [15:0] Tile_X03_Y00_io2f_16;
	// wire [8:0] Tile_X03_Y00_hi;
	// wire [7:0] Tile_X03_Y00_lo;
	// wire [0:0] Tile_X03_Y01_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y01_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y01_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y01_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y01_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y01_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y01_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y01_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y01_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y01_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y01_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y01_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X03_Y01_clk_out;
	// wire Tile_X03_Y01_clk_pass_through_out_bot;
	// wire [31:0] Tile_X03_Y01_config_out_config_addr;
	// wire [31:0] Tile_X03_Y01_config_out_config_data;
	// wire [0:0] Tile_X03_Y01_config_out_read;
	// wire [0:0] Tile_X03_Y01_config_out_write;
	// wire [8:0] Tile_X03_Y01_hi_unq1;
	// wire [7:0] Tile_X03_Y01_lo_unq1;
	// wire [31:0] Tile_X03_Y01_read_config_data;
	// wire Tile_X03_Y01_reset_out;
	// wire [0:0] Tile_X03_Y01_stall_out;
	// wire [8:0] Tile_X03_Y01_hi_out;
	// wire [7:0] Tile_X03_Y01_lo_out;
	// wire [15:0] Tile_X03_Y01_tile_id_in;
	// wire [0:0] Tile_X03_Y02_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y02_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y02_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y02_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y02_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y02_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y02_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y02_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y02_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y02_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y02_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y02_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X03_Y02_clk_out;
	// wire Tile_X03_Y02_clk_pass_through_out_bot;
	// wire [31:0] Tile_X03_Y02_config_out_config_addr;
	// wire [31:0] Tile_X03_Y02_config_out_config_data;
	// wire [0:0] Tile_X03_Y02_config_out_read;
	// wire [0:0] Tile_X03_Y02_config_out_write;
	// wire [8:0] Tile_X03_Y02_hi_unq1;
	// wire [7:0] Tile_X03_Y02_lo_unq1;
	// wire [31:0] Tile_X03_Y02_read_config_data;
	// wire Tile_X03_Y02_reset_out;
	// wire [0:0] Tile_X03_Y02_stall_out;
	// wire [8:0] Tile_X03_Y02_hi_out;
	// wire [7:0] Tile_X03_Y02_lo_out;
	// wire [15:0] Tile_X03_Y02_tile_id_in;
	// wire [0:0] Tile_X03_Y03_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y03_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y03_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y03_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y03_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y03_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y03_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y03_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y03_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y03_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y03_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y03_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X03_Y03_clk_out;
	// wire Tile_X03_Y03_clk_pass_through_out_bot;
	// wire [31:0] Tile_X03_Y03_config_out_config_addr;
	// wire [31:0] Tile_X03_Y03_config_out_config_data;
	// wire [0:0] Tile_X03_Y03_config_out_read;
	// wire [0:0] Tile_X03_Y03_config_out_write;
	// wire [8:0] Tile_X03_Y03_hi_unq1;
	// wire [7:0] Tile_X03_Y03_lo_unq1;
	// wire [31:0] Tile_X03_Y03_read_config_data;
	// wire Tile_X03_Y03_reset_out;
	// wire [0:0] Tile_X03_Y03_stall_out;
	// wire [8:0] Tile_X03_Y03_hi_out;
	// wire [7:0] Tile_X03_Y03_lo_out;
	// wire [15:0] Tile_X03_Y03_tile_id_in;
	// wire [0:0] Tile_X03_Y04_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y04_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y04_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y04_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y04_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y04_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y04_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y04_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y04_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y04_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y04_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y04_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X03_Y04_clk_out;
	// wire Tile_X03_Y04_clk_pass_through_out_bot;
	// wire [31:0] Tile_X03_Y04_config_out_config_addr;
	// wire [31:0] Tile_X03_Y04_config_out_config_data;
	// wire [0:0] Tile_X03_Y04_config_out_read;
	// wire [0:0] Tile_X03_Y04_config_out_write;
	// wire [8:0] Tile_X03_Y04_hi_unq1;
	// wire [7:0] Tile_X03_Y04_lo_unq1;
	// wire [31:0] Tile_X03_Y04_read_config_data;
	// wire Tile_X03_Y04_reset_out;
	// wire [0:0] Tile_X03_Y04_stall_out;
	// wire [8:0] Tile_X03_Y04_hi_out;
	// wire [7:0] Tile_X03_Y04_lo_out;
	// wire [15:0] Tile_X03_Y04_tile_id_in;
	// wire [0:0] Tile_X03_Y05_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y05_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y05_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y05_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y05_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y05_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y05_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y05_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y05_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y05_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y05_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y05_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y05_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y05_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y05_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y05_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y05_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y05_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y05_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y05_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y05_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y05_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y05_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y05_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X03_Y05_clk_out;
	// wire Tile_X03_Y05_clk_pass_through_out_bot;
	// wire [31:0] Tile_X03_Y05_config_out_config_addr;
	// wire [31:0] Tile_X03_Y05_config_out_config_data;
	// wire [0:0] Tile_X03_Y05_config_out_read;
	// wire [0:0] Tile_X03_Y05_config_out_write;
	// wire [8:0] Tile_X03_Y05_hi_unq1;
	// wire [7:0] Tile_X03_Y05_lo_unq1;
	// wire [31:0] Tile_X03_Y05_read_config_data;
	// wire Tile_X03_Y05_reset_out;
	// wire [0:0] Tile_X03_Y05_stall_out;
	// wire [8:0] Tile_X03_Y05_hi_out;
	// wire [7:0] Tile_X03_Y05_lo_out;
	// wire [15:0] Tile_X03_Y05_tile_id_in;
	// wire [0:0] Tile_X03_Y06_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y06_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y06_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y06_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y06_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y06_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y06_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y06_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y06_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y06_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y06_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y06_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y06_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y06_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y06_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y06_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y06_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y06_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y06_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y06_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y06_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y06_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y06_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y06_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X03_Y06_clk_out;
	// wire Tile_X03_Y06_clk_pass_through_out_bot;
	// wire [31:0] Tile_X03_Y06_config_out_config_addr;
	// wire [31:0] Tile_X03_Y06_config_out_config_data;
	// wire [0:0] Tile_X03_Y06_config_out_read;
	// wire [0:0] Tile_X03_Y06_config_out_write;
	// wire [8:0] Tile_X03_Y06_hi_unq1;
	// wire [7:0] Tile_X03_Y06_lo_unq1;
	// wire [31:0] Tile_X03_Y06_read_config_data;
	// wire Tile_X03_Y06_reset_out;
	// wire [0:0] Tile_X03_Y06_stall_out;
	// wire [8:0] Tile_X03_Y06_hi_out;
	// wire [7:0] Tile_X03_Y06_lo_out;
	// wire [15:0] Tile_X03_Y06_tile_id_in;
	// wire [0:0] Tile_X03_Y07_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y07_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y07_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y07_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y07_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y07_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y07_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y07_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y07_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y07_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y07_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y07_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y07_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y07_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y07_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y07_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y07_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y07_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y07_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y07_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y07_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y07_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y07_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y07_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X03_Y07_clk_out;
	// wire Tile_X03_Y07_clk_pass_through_out_bot;
	// wire [31:0] Tile_X03_Y07_config_out_config_addr;
	// wire [31:0] Tile_X03_Y07_config_out_config_data;
	// wire [0:0] Tile_X03_Y07_config_out_read;
	// wire [0:0] Tile_X03_Y07_config_out_write;
	// wire [8:0] Tile_X03_Y07_hi_unq1;
	// wire [7:0] Tile_X03_Y07_lo_unq1;
	// wire [31:0] Tile_X03_Y07_read_config_data;
	// wire Tile_X03_Y07_reset_out;
	// wire [0:0] Tile_X03_Y07_stall_out;
	// wire [8:0] Tile_X03_Y07_hi_out;
	// wire [7:0] Tile_X03_Y07_lo_out;
	// wire [15:0] Tile_X03_Y07_tile_id_in;
	// wire [0:0] Tile_X03_Y08_SB_T0_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y08_SB_T0_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y08_SB_T0_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y08_SB_T0_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y08_SB_T0_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y08_SB_T0_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y08_SB_T0_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y08_SB_T0_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y08_SB_T1_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y08_SB_T1_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y08_SB_T1_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y08_SB_T1_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y08_SB_T1_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y08_SB_T1_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y08_SB_T1_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y08_SB_T1_WEST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y08_SB_T2_EAST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y08_SB_T2_EAST_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y08_SB_T2_NORTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y08_SB_T2_NORTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y08_SB_T2_SOUTH_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y08_SB_T2_SOUTH_SB_OUT_B16;
	// wire [0:0] Tile_X03_Y08_SB_T2_WEST_SB_OUT_B1;
	// wire [15:0] Tile_X03_Y08_SB_T2_WEST_SB_OUT_B16;
	// wire Tile_X03_Y08_clk_out;
	// wire Tile_X03_Y08_clk_pass_through_out_bot;
	// wire [31:0] Tile_X03_Y08_config_out_config_addr;
	// wire [31:0] Tile_X03_Y08_config_out_config_data;
	// wire [0:0] Tile_X03_Y08_config_out_read;
	// wire [0:0] Tile_X03_Y08_config_out_write;
	// wire [8:0] Tile_X03_Y08_hi_unq1;
	// wire [7:0] Tile_X03_Y08_lo_unq1;
	// wire [31:0] Tile_X03_Y08_read_config_data;
	// wire Tile_X03_Y08_reset_out;
	// wire [0:0] Tile_X03_Y08_stall_out;
	// wire [8:0] Tile_X03_Y08_hi_out;
	// wire [7:0] Tile_X03_Y08_lo_out;
	// wire [15:0] Tile_X03_Y08_tile_id_in;
	wire [0:0] const_0_1_out;
	wire [15:0] const_0_16_out;
	wire [31:0] const_0_32_out;
	wire [31:0] read_config_data_or_final_O;
	wire [15:0] Tile_X00_Y00_tile_id;
	assign Tile_X00_Y00_tile_id = {Tile_X00_Y00_lo[7], Tile_X00_Y00_lo[7:6], Tile_X00_Y00_lo[6:5], Tile_X00_Y00_lo[5:4], Tile_X00_Y00_lo[4:3], Tile_X00_Y00_lo[3:2], Tile_X00_Y00_lo[2:1], Tile_X00_Y00_lo[1:0], Tile_X00_Y00_lo[0]};
	Tile_io_core Tile_X00_Y00(
		.tile_id(Tile_X00_Y00_tile_id),
		.glb2io_1(glb2io_1_X00_Y00),
		.f2io_1(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B1),
		.io2glb_1(Tile_X00_Y00_io2glb_1),
		.io2f_1(Tile_X00_Y00_io2f_1),
		.glb2io_16(glb2io_16_X00_Y00),
		.f2io_16(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B16),
		.io2glb_16(Tile_X00_Y00_io2glb_16),
		.io2f_16(Tile_X00_Y00_io2f_16),
		.hi(Tile_X00_Y00_hi),
		.lo(Tile_X00_Y00_lo)
	);
	Tile_MemCore Tile_X00_Y01(
		.SB_T0_EAST_SB_IN_B1(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_EAST_SB_IN_B16(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B16),
		.SB_T0_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B16(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B16),
		.SB_T0_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
		.SB_T0_NORTH_SB_IN_B16(Tile_X00_Y00_io2f_16),
		.SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B16),
		.SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B16),
		.SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B16),
		.SB_T0_WEST_SB_IN_B1(const_0_1_out),
		.SB_T0_WEST_SB_IN_B16(const_0_16_out),
		.SB_T0_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B16(Tile_X00_Y01_SB_T0_WEST_SB_OUT_B16),
		.SB_T1_EAST_SB_IN_B1(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_EAST_SB_IN_B16(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B16),
		.SB_T1_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B16(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B16),
		.SB_T1_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
		.SB_T1_NORTH_SB_IN_B16(Tile_X00_Y00_io2f_16),
		.SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B16),
		.SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B16),
		.SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B16),
		.SB_T1_WEST_SB_IN_B1(const_0_1_out),
		.SB_T1_WEST_SB_IN_B16(const_0_16_out),
		.SB_T1_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B16(Tile_X00_Y01_SB_T1_WEST_SB_OUT_B16),
		.SB_T2_EAST_SB_IN_B1(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_EAST_SB_IN_B16(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B16),
		.SB_T2_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B16(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B16),
		.SB_T2_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
		.SB_T2_NORTH_SB_IN_B16(Tile_X00_Y00_io2f_16),
		.SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B16),
		.SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B16),
		.SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B16),
		.SB_T2_WEST_SB_IN_B1(const_0_1_out),
		.SB_T2_WEST_SB_IN_B16(const_0_16_out),
		.SB_T2_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B16(Tile_X00_Y01_SB_T2_WEST_SB_OUT_B16),
		.clk(clk),
		.clk_out(Tile_X00_Y01_clk_out),
		.clk_pass_through(clk),
		.clk_pass_through_out_bot(Tile_X00_Y01_clk_pass_through_out_bot),
		.config_config_addr(config_0_config_addr),
		.config_config_data(config_0_config_data),
		.config_out_config_addr(Tile_X00_Y01_config_out_config_addr),
		.config_out_config_data(Tile_X00_Y01_config_out_config_data),
		.config_out_read(Tile_X00_Y01_config_out_read),
		.config_out_write(Tile_X00_Y01_config_out_write),
		.config_read(config_0_read),
		.config_write(config_0_write),
		.hi(Tile_X00_Y01_hi),
		.lo(Tile_X00_Y01_lo_unq1),
		.read_config_data(Tile_X00_Y01_read_config_data),
		.read_config_data_in(const_0_32_out),
		.reset(reset),
		.reset_out(Tile_X00_Y01_reset_out),
		.stall(stall[0]),
		.stall_out(Tile_X00_Y01_stall_out),
		.tile_id(Tile_X00_Y01_tile_id_in)
	);
	mantle_wire__typeBit8 Tile_X00_Y01_lo(
		.in(Tile_X00_Y01_lo_unq1),
		.out(Tile_X00_Y01_lo_out)
	);
	wire [15:0] Tile_X00_Y01_tile_id_out;
	assign Tile_X00_Y01_tile_id_out = {Tile_X00_Y01_lo_out[7], Tile_X00_Y01_lo_out[7:6], Tile_X00_Y01_lo_out[6:5], Tile_X00_Y01_lo_out[5:4], Tile_X00_Y01_lo_out[4:3], Tile_X00_Y01_lo_out[3:2], Tile_X00_Y01_lo_out[2:1], Tile_X00_Y01_lo_out[1:0], Tile_X00_Y01_hi[0]};
	mantle_wire__typeBitIn16 Tile_X00_Y01_tile_id(
		.in(Tile_X00_Y01_tile_id_in),
		.out(Tile_X00_Y01_tile_id_out)
	);
	Tile_PE Tile_X00_Y02(
		.SB_T0_EAST_SB_IN_B1(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_EAST_SB_IN_B16(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B16),
		.SB_T0_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B16(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B16),
		.SB_T0_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_IN_B16(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B16),
		.SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B16),
		// .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B1),
		// .SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B16),
		.SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B16),
		.SB_T0_WEST_SB_IN_B1(const_0_1_out),
		.SB_T0_WEST_SB_IN_B16(const_0_16_out),
		.SB_T0_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B16(Tile_X00_Y02_SB_T0_WEST_SB_OUT_B16),
		.SB_T1_EAST_SB_IN_B1(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_EAST_SB_IN_B16(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B16),
		.SB_T1_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B16(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B16),
		.SB_T1_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_IN_B16(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B16),
		.SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B16),
		// .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B1),
		// .SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B16),
		.SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B16),
		.SB_T1_WEST_SB_IN_B1(const_0_1_out),
		.SB_T1_WEST_SB_IN_B16(const_0_16_out),
		.SB_T1_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B16(Tile_X00_Y02_SB_T1_WEST_SB_OUT_B16),
		.SB_T2_EAST_SB_IN_B1(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_EAST_SB_IN_B16(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B16),
		.SB_T2_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B16(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B16),
		.SB_T2_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_IN_B16(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B16),
		.SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B16),
		// .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B1),
		// .SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B16),
		.SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B16),
		.SB_T2_WEST_SB_IN_B1(const_0_1_out),
		.SB_T2_WEST_SB_IN_B16(const_0_16_out),
		.SB_T2_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B16(Tile_X00_Y02_SB_T2_WEST_SB_OUT_B16),
		.clk(Tile_X00_Y01_clk_out),
		.clk_out(Tile_X00_Y02_clk_out),
		.clk_pass_through(Tile_X00_Y01_clk_pass_through_out_bot),
		.clk_pass_through_out_bot(Tile_X00_Y02_clk_pass_through_out_bot),
		.config_config_addr(Tile_X00_Y01_config_out_config_addr),
		.config_config_data(Tile_X00_Y01_config_out_config_data),
		.config_out_config_addr(Tile_X00_Y02_config_out_config_addr),
		.config_out_config_data(Tile_X00_Y02_config_out_config_data),
		.config_out_read(Tile_X00_Y02_config_out_read),
		.config_out_write(Tile_X00_Y02_config_out_write),
		.config_read(Tile_X00_Y01_config_out_read),
		.config_write(Tile_X00_Y01_config_out_write),
		.hi(Tile_X00_Y02_hi),
		.lo(Tile_X00_Y02_lo_unq1),
		.read_config_data(Tile_X00_Y02_read_config_data),
		.read_config_data_in(Tile_X00_Y01_read_config_data),
		.reset(Tile_X00_Y01_reset_out),
		.reset_out(Tile_X00_Y02_reset_out),
		.stall(Tile_X00_Y01_stall_out),
		.stall_out(Tile_X00_Y02_stall_out),
		.tile_id(Tile_X00_Y02_tile_id_in)
	);
	mantle_wire__typeBit8 Tile_X00_Y02_lo(
		.in(Tile_X00_Y02_lo_unq1),
		.out(Tile_X00_Y02_lo_out)
	);
	wire [15:0] Tile_X00_Y02_tile_id_out;
	assign Tile_X00_Y02_tile_id_out = {Tile_X00_Y02_lo_out[7], Tile_X00_Y02_lo_out[7:6], Tile_X00_Y02_lo_out[6:5], Tile_X00_Y02_lo_out[5:4], Tile_X00_Y02_lo_out[4:3], Tile_X00_Y02_lo_out[3:2], Tile_X00_Y02_lo_out[2:1], Tile_X00_Y02_lo_out[1], Tile_X00_Y02_hi[1], Tile_X00_Y02_lo_out[0]};
	mantle_wire__typeBitIn16 Tile_X00_Y02_tile_id(
		.in(Tile_X00_Y02_tile_id_in),
		.out(Tile_X00_Y02_tile_id_out)
	);
	// Tile_PE Tile_X00_Y03(
	// 	.SB_T0_EAST_SB_IN_B1(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_IN_B16(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(const_0_1_out),
	// 	.SB_T0_WEST_SB_IN_B16(const_0_16_out),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X00_Y03_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_IN_B16(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(const_0_1_out),
	// 	.SB_T1_WEST_SB_IN_B16(const_0_16_out),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X00_Y03_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_IN_B16(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(const_0_1_out),
	// 	.SB_T2_WEST_SB_IN_B16(const_0_16_out),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X00_Y03_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X00_Y02_clk_out),
	// 	.clk_out(Tile_X00_Y03_clk_out),
	// 	.clk_pass_through(Tile_X00_Y02_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X00_Y03_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X00_Y02_config_out_config_addr),
	// 	.config_config_data(Tile_X00_Y02_config_out_config_data),
	// 	.config_out_config_addr(Tile_X00_Y03_config_out_config_addr),
	// 	.config_out_config_data(Tile_X00_Y03_config_out_config_data),
	// 	.config_out_read(Tile_X00_Y03_config_out_read),
	// 	.config_out_write(Tile_X00_Y03_config_out_write),
	// 	.config_read(Tile_X00_Y02_config_out_read),
	// 	.config_write(Tile_X00_Y02_config_out_write),
	// 	.hi(Tile_X00_Y03_hi_unq1),
	// 	.lo(Tile_X00_Y03_lo_unq1),
	// 	.read_config_data(Tile_X00_Y03_read_config_data),
	// 	.read_config_data_in(Tile_X00_Y02_read_config_data),
	// 	.reset(Tile_X00_Y02_reset_out),
	// 	.reset_out(Tile_X00_Y03_reset_out),
	// 	.stall(Tile_X00_Y02_stall_out),
	// 	.stall_out(Tile_X00_Y03_stall_out),
	// 	.tile_id(Tile_X00_Y03_tile_id_in)
	// );
	// mantle_wire__typeBit9 Tile_X00_Y03_hi(
	// 	.in(Tile_X00_Y03_hi_unq1),
	// 	.out(Tile_X00_Y03_hi_out)
	// );
	// mantle_wire__typeBit8 Tile_X00_Y03_lo(
	// 	.in(Tile_X00_Y03_lo_unq1),
	// 	.out(Tile_X00_Y03_lo_out)
	// );
	// wire [15:0] Tile_X00_Y03_tile_id_out;
	// assign Tile_X00_Y03_tile_id_out = {Tile_X00_Y03_lo_out[7], Tile_X00_Y03_lo_out[7:6], Tile_X00_Y03_lo_out[6:5], Tile_X00_Y03_lo_out[5:4], Tile_X00_Y03_lo_out[4:3], Tile_X00_Y03_lo_out[3:2], Tile_X00_Y03_lo_out[2:1], Tile_X00_Y03_lo_out[1], Tile_X00_Y03_hi_out[1:0]};
	// mantle_wire__typeBitIn16 Tile_X00_Y03_tile_id(
	// 	.in(Tile_X00_Y03_tile_id_in),
	// 	.out(Tile_X00_Y03_tile_id_out)
	// );
	// Tile_PE Tile_X00_Y04(
	// 	.SB_T0_EAST_SB_IN_B1(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_IN_B16(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y05_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y05_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(const_0_1_out),
	// 	.SB_T0_WEST_SB_IN_B16(const_0_16_out),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X00_Y04_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_IN_B16(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y05_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y05_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(const_0_1_out),
	// 	.SB_T1_WEST_SB_IN_B16(const_0_16_out),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X00_Y04_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_IN_B16(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y05_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y05_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(const_0_1_out),
	// 	.SB_T2_WEST_SB_IN_B16(const_0_16_out),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X00_Y04_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X00_Y03_clk_out),
	// 	.clk_out(Tile_X00_Y04_clk_out),
	// 	.clk_pass_through(Tile_X00_Y03_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X00_Y04_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X00_Y03_config_out_config_addr),
	// 	.config_config_data(Tile_X00_Y03_config_out_config_data),
	// 	.config_out_config_addr(Tile_X00_Y04_config_out_config_addr),
	// 	.config_out_config_data(Tile_X00_Y04_config_out_config_data),
	// 	.config_out_read(Tile_X00_Y04_config_out_read),
	// 	.config_out_write(Tile_X00_Y04_config_out_write),
	// 	.config_read(Tile_X00_Y03_config_out_read),
	// 	.config_write(Tile_X00_Y03_config_out_write),
	// 	.hi(Tile_X00_Y04_hi),
	// 	.lo(Tile_X00_Y04_lo_unq1),
	// 	.read_config_data(Tile_X00_Y04_read_config_data),
	// 	.read_config_data_in(Tile_X00_Y03_read_config_data),
	// 	.reset(Tile_X00_Y03_reset_out),
	// 	.reset_out(Tile_X00_Y04_reset_out),
	// 	.stall(Tile_X00_Y03_stall_out),
	// 	.stall_out(Tile_X00_Y04_stall_out),
	// 	.tile_id(Tile_X00_Y04_tile_id_in)
	// );
	// mantle_wire__typeBit8 Tile_X00_Y04_lo(
	// 	.in(Tile_X00_Y04_lo_unq1),
	// 	.out(Tile_X00_Y04_lo_out)
	// );
	// wire [15:0] Tile_X00_Y04_tile_id_out;
	// assign Tile_X00_Y04_tile_id_out = {Tile_X00_Y04_lo_out[7], Tile_X00_Y04_lo_out[7:6], Tile_X00_Y04_lo_out[6:5], Tile_X00_Y04_lo_out[5:4], Tile_X00_Y04_lo_out[4:3], Tile_X00_Y04_lo_out[3:2], Tile_X00_Y04_lo_out[2:1], Tile_X00_Y04_hi[1], Tile_X00_Y04_lo_out[0], Tile_X00_Y04_lo_out[0]};
	// mantle_wire__typeBitIn16 Tile_X00_Y04_tile_id(
	// 	.in(Tile_X00_Y04_tile_id_in),
	// 	.out(Tile_X00_Y04_tile_id_out)
	// );
	// Tile_MemCore Tile_X00_Y05(
	// 	.SB_T0_EAST_SB_IN_B1(Tile_X01_Y05_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_IN_B16(Tile_X01_Y05_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X00_Y05_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X00_Y05_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y05_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y05_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y06_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y06_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y05_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y05_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(const_0_1_out),
	// 	.SB_T0_WEST_SB_IN_B16(const_0_16_out),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X00_Y05_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X00_Y05_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(Tile_X01_Y05_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_IN_B16(Tile_X01_Y05_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X00_Y05_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X00_Y05_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y05_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y05_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y06_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y06_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y05_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y05_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(const_0_1_out),
	// 	.SB_T1_WEST_SB_IN_B16(const_0_16_out),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X00_Y05_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X00_Y05_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(Tile_X01_Y05_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_IN_B16(Tile_X01_Y05_SB_T2_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X00_Y05_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X00_Y05_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y05_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y05_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y06_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y06_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y05_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y05_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(const_0_1_out),
	// 	.SB_T2_WEST_SB_IN_B16(const_0_16_out),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X00_Y05_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X00_Y05_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X00_Y04_clk_out),
	// 	.clk_out(Tile_X00_Y05_clk_out),
	// 	.clk_pass_through(Tile_X00_Y04_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X00_Y05_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X00_Y04_config_out_config_addr),
	// 	.config_config_data(Tile_X00_Y04_config_out_config_data),
	// 	.config_out_config_addr(Tile_X00_Y05_config_out_config_addr),
	// 	.config_out_config_data(Tile_X00_Y05_config_out_config_data),
	// 	.config_out_read(Tile_X00_Y05_config_out_read),
	// 	.config_out_write(Tile_X00_Y05_config_out_write),
	// 	.config_read(Tile_X00_Y04_config_out_read),
	// 	.config_write(Tile_X00_Y04_config_out_write),
	// 	.hi(Tile_X00_Y05_hi),
	// 	.lo(Tile_X00_Y05_lo_unq1),
	// 	.read_config_data(Tile_X00_Y05_read_config_data),
	// 	.read_config_data_in(Tile_X00_Y04_read_config_data),
	// 	.reset(Tile_X00_Y04_reset_out),
	// 	.reset_out(Tile_X00_Y05_reset_out),
	// 	.stall(Tile_X00_Y04_stall_out),
	// 	.stall_out(Tile_X00_Y05_stall_out),
	// 	.tile_id(Tile_X00_Y05_tile_id_in)
	// );
	// mantle_wire__typeBit8 Tile_X00_Y05_lo(
	// 	.in(Tile_X00_Y05_lo_unq1),
	// 	.out(Tile_X00_Y05_lo_out)
	// );
	// wire [15:0] Tile_X00_Y05_tile_id_out;
	// assign Tile_X00_Y05_tile_id_out = {Tile_X00_Y05_lo_out[7], Tile_X00_Y05_lo_out[7:6], Tile_X00_Y05_lo_out[6:5], Tile_X00_Y05_lo_out[5:4], Tile_X00_Y05_lo_out[4:3], Tile_X00_Y05_lo_out[3:2], Tile_X00_Y05_lo_out[2:1], Tile_X00_Y05_hi[1], Tile_X00_Y05_lo_out[0], Tile_X00_Y05_hi[0]};
	// mantle_wire__typeBitIn16 Tile_X00_Y05_tile_id(
	// 	.in(Tile_X00_Y05_tile_id_in),
	// 	.out(Tile_X00_Y05_tile_id_out)
	// );
	// Tile_PE Tile_X00_Y06(
	// 	.SB_T0_EAST_SB_IN_B1(Tile_X01_Y06_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_IN_B16(Tile_X01_Y06_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X00_Y06_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X00_Y06_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X00_Y05_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X00_Y05_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y06_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y06_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y07_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y07_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y06_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y06_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(const_0_1_out),
	// 	.SB_T0_WEST_SB_IN_B16(const_0_16_out),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X00_Y06_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X00_Y06_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(Tile_X01_Y06_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_IN_B16(Tile_X01_Y06_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X00_Y06_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X00_Y06_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X00_Y05_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X00_Y05_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y06_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y06_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y07_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y07_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y06_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y06_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(const_0_1_out),
	// 	.SB_T1_WEST_SB_IN_B16(const_0_16_out),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X00_Y06_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X00_Y06_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(Tile_X01_Y06_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_IN_B16(Tile_X01_Y06_SB_T2_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X00_Y06_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X00_Y06_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X00_Y05_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X00_Y05_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y06_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y06_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y07_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y07_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y06_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y06_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(const_0_1_out),
	// 	.SB_T2_WEST_SB_IN_B16(const_0_16_out),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X00_Y06_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X00_Y06_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X00_Y05_clk_out),
	// 	.clk_out(Tile_X00_Y06_clk_out),
	// 	.clk_pass_through(Tile_X00_Y05_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X00_Y06_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X00_Y05_config_out_config_addr),
	// 	.config_config_data(Tile_X00_Y05_config_out_config_data),
	// 	.config_out_config_addr(Tile_X00_Y06_config_out_config_addr),
	// 	.config_out_config_data(Tile_X00_Y06_config_out_config_data),
	// 	.config_out_read(Tile_X00_Y06_config_out_read),
	// 	.config_out_write(Tile_X00_Y06_config_out_write),
	// 	.config_read(Tile_X00_Y05_config_out_read),
	// 	.config_write(Tile_X00_Y05_config_out_write),
	// 	.hi(Tile_X00_Y06_hi),
	// 	.lo(Tile_X00_Y06_lo_unq1),
	// 	.read_config_data(Tile_X00_Y06_read_config_data),
	// 	.read_config_data_in(Tile_X00_Y05_read_config_data),
	// 	.reset(Tile_X00_Y05_reset_out),
	// 	.reset_out(Tile_X00_Y06_reset_out),
	// 	.stall(Tile_X00_Y05_stall_out),
	// 	.stall_out(Tile_X00_Y06_stall_out),
	// 	.tile_id(Tile_X00_Y06_tile_id_in)
	// );
	// mantle_wire__typeBit8 Tile_X00_Y06_lo(
	// 	.in(Tile_X00_Y06_lo_unq1),
	// 	.out(Tile_X00_Y06_lo_out)
	// );
	// wire [15:0] Tile_X00_Y06_tile_id_out;
	// assign Tile_X00_Y06_tile_id_out = {Tile_X00_Y06_lo_out[7], Tile_X00_Y06_lo_out[7:6], Tile_X00_Y06_lo_out[6:5], Tile_X00_Y06_lo_out[5:4], Tile_X00_Y06_lo_out[4:3], Tile_X00_Y06_lo_out[3:2], Tile_X00_Y06_lo_out[2:1], Tile_X00_Y06_hi[1], Tile_X00_Y06_hi[1], Tile_X00_Y06_lo_out[0]};
	// mantle_wire__typeBitIn16 Tile_X00_Y06_tile_id(
	// 	.in(Tile_X00_Y06_tile_id_in),
	// 	.out(Tile_X00_Y06_tile_id_out)
	// );
	// Tile_PE Tile_X00_Y07(
	// 	.SB_T0_EAST_SB_IN_B1(Tile_X01_Y07_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_IN_B16(Tile_X01_Y07_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X00_Y07_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X00_Y07_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X00_Y06_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X00_Y06_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y07_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y07_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y08_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y08_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y07_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y07_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(const_0_1_out),
	// 	.SB_T0_WEST_SB_IN_B16(const_0_16_out),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X00_Y07_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X00_Y07_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(Tile_X01_Y07_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_IN_B16(Tile_X01_Y07_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X00_Y07_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X00_Y07_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X00_Y06_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X00_Y06_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y07_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y07_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y08_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y08_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y07_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y07_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(const_0_1_out),
	// 	.SB_T1_WEST_SB_IN_B16(const_0_16_out),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X00_Y07_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X00_Y07_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(Tile_X01_Y07_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_IN_B16(Tile_X01_Y07_SB_T2_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X00_Y07_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X00_Y07_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X00_Y06_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X00_Y06_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y07_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y07_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y08_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y08_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y07_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y07_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(const_0_1_out),
	// 	.SB_T2_WEST_SB_IN_B16(const_0_16_out),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X00_Y07_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X00_Y07_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X00_Y06_clk_out),
	// 	.clk_out(Tile_X00_Y07_clk_out),
	// 	.clk_pass_through(Tile_X00_Y06_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X00_Y07_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X00_Y06_config_out_config_addr),
	// 	.config_config_data(Tile_X00_Y06_config_out_config_data),
	// 	.config_out_config_addr(Tile_X00_Y07_config_out_config_addr),
	// 	.config_out_config_data(Tile_X00_Y07_config_out_config_data),
	// 	.config_out_read(Tile_X00_Y07_config_out_read),
	// 	.config_out_write(Tile_X00_Y07_config_out_write),
	// 	.config_read(Tile_X00_Y06_config_out_read),
	// 	.config_write(Tile_X00_Y06_config_out_write),
	// 	.hi(Tile_X00_Y07_hi_unq1),
	// 	.lo(Tile_X00_Y07_lo_unq1),
	// 	.read_config_data(Tile_X00_Y07_read_config_data),
	// 	.read_config_data_in(Tile_X00_Y06_read_config_data),
	// 	.reset(Tile_X00_Y06_reset_out),
	// 	.reset_out(Tile_X00_Y07_reset_out),
	// 	.stall(Tile_X00_Y06_stall_out),
	// 	.stall_out(Tile_X00_Y07_stall_out),
	// 	.tile_id(Tile_X00_Y07_tile_id_in)
	// );
	// mantle_wire__typeBit9 Tile_X00_Y07_hi(
	// 	.in(Tile_X00_Y07_hi_unq1),
	// 	.out(Tile_X00_Y07_hi_out)
	// );
	// mantle_wire__typeBit8 Tile_X00_Y07_lo(
	// 	.in(Tile_X00_Y07_lo_unq1),
	// 	.out(Tile_X00_Y07_lo_out)
	// );
	// wire [15:0] Tile_X00_Y07_tile_id_out;
	// assign Tile_X00_Y07_tile_id_out = {Tile_X00_Y07_lo_out[7], Tile_X00_Y07_lo_out[7:6], Tile_X00_Y07_lo_out[6:5], Tile_X00_Y07_lo_out[5:4], Tile_X00_Y07_lo_out[4:3], Tile_X00_Y07_lo_out[3:2], Tile_X00_Y07_lo_out[2:1], Tile_X00_Y07_hi_out[1], Tile_X00_Y07_hi_out[1:0]};
	// mantle_wire__typeBitIn16 Tile_X00_Y07_tile_id(
	// 	.in(Tile_X00_Y07_tile_id_in),
	// 	.out(Tile_X00_Y07_tile_id_out)
	// );
	// Tile_PE Tile_X00_Y08(
	// 	.SB_T0_EAST_SB_IN_B1(Tile_X01_Y08_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_IN_B16(Tile_X01_Y08_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X00_Y08_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X00_Y08_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X00_Y07_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X00_Y07_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y08_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y08_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
	// 	.SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y08_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y08_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(const_0_1_out),
	// 	.SB_T0_WEST_SB_IN_B16(const_0_16_out),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X00_Y08_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X00_Y08_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(Tile_X01_Y08_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_IN_B16(Tile_X01_Y08_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X00_Y08_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X00_Y08_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X00_Y07_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X00_Y07_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y08_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y08_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
	// 	.SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y08_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y08_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(const_0_1_out),
	// 	.SB_T1_WEST_SB_IN_B16(const_0_16_out),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X00_Y08_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X00_Y08_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(Tile_X01_Y08_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_IN_B16(Tile_X01_Y08_SB_T2_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X00_Y08_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X00_Y08_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X00_Y07_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X00_Y07_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y08_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y08_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
	// 	.SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y08_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y08_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(const_0_1_out),
	// 	.SB_T2_WEST_SB_IN_B16(const_0_16_out),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X00_Y08_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X00_Y08_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X00_Y07_clk_out),
	// 	.clk_out(Tile_X00_Y08_clk_out),
	// 	.clk_pass_through(Tile_X00_Y07_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X00_Y08_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X00_Y07_config_out_config_addr),
	// 	.config_config_data(Tile_X00_Y07_config_out_config_data),
	// 	.config_out_config_addr(Tile_X00_Y08_config_out_config_addr),
	// 	.config_out_config_data(Tile_X00_Y08_config_out_config_data),
	// 	.config_out_read(Tile_X00_Y08_config_out_read),
	// 	.config_out_write(Tile_X00_Y08_config_out_write),
	// 	.config_read(Tile_X00_Y07_config_out_read),
	// 	.config_write(Tile_X00_Y07_config_out_write),
	// 	.hi(Tile_X00_Y08_hi),
	// 	.lo(Tile_X00_Y08_lo_unq1),
	// 	.read_config_data(Tile_X00_Y08_read_config_data),
	// 	.read_config_data_in(Tile_X00_Y07_read_config_data),
	// 	.reset(Tile_X00_Y07_reset_out),
	// 	.reset_out(Tile_X00_Y08_reset_out),
	// 	.stall(Tile_X00_Y07_stall_out),
	// 	.stall_out(Tile_X00_Y08_stall_out),
	// 	.tile_id(Tile_X00_Y08_tile_id_in)
	// );
	// mantle_wire__typeBit8 Tile_X00_Y08_lo(
	// 	.in(Tile_X00_Y08_lo_unq1),
	// 	.out(Tile_X00_Y08_lo_out)
	// );
	// wire [15:0] Tile_X00_Y08_tile_id_out;
	// assign Tile_X00_Y08_tile_id_out = {Tile_X00_Y08_lo_out[7], Tile_X00_Y08_lo_out[7:6], Tile_X00_Y08_lo_out[6:5], Tile_X00_Y08_lo_out[5:4], Tile_X00_Y08_lo_out[4:3], Tile_X00_Y08_lo_out[3:2], Tile_X00_Y08_lo_out[2], Tile_X00_Y08_hi[2], Tile_X00_Y08_lo_out[1:0], Tile_X00_Y08_lo_out[0]};
	// mantle_wire__typeBitIn16 Tile_X00_Y08_tile_id(
	// 	.in(Tile_X00_Y08_tile_id_in),
	// 	.out(Tile_X00_Y08_tile_id_out)
	// );
	wire [15:0] Tile_X01_Y00_tile_id;
	assign Tile_X01_Y00_tile_id = {Tile_X01_Y00_lo[7], Tile_X01_Y00_lo[7:6], Tile_X01_Y00_lo[6:5], Tile_X01_Y00_lo[5:4], Tile_X01_Y00_hi[4], Tile_X01_Y00_lo[3], Tile_X01_Y00_lo[3:2], Tile_X01_Y00_lo[2:1], Tile_X01_Y00_lo[1:0], Tile_X01_Y00_lo[0]};
	Tile_io_core Tile_X01_Y00(
		.tile_id(Tile_X01_Y00_tile_id),
		.glb2io_1(glb2io_1_X01_Y00),
		.f2io_1(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B1),
		.io2glb_1(Tile_X01_Y00_io2glb_1),
		.io2f_1(Tile_X01_Y00_io2f_1),
		.glb2io_16(glb2io_16_X01_Y00),
		.f2io_16(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B16),
		.io2glb_16(Tile_X01_Y00_io2glb_16),
		.io2f_16(Tile_X01_Y00_io2f_16),
		.hi(Tile_X01_Y00_hi),
		.lo(Tile_X01_Y00_lo)
	);
	Tile_MemCore Tile_X01_Y01(
		// .SB_T0_EAST_SB_IN_B1(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B1),
		// .SB_T0_EAST_SB_IN_B16(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B16),
		.SB_T0_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B16(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B16),
		.SB_T0_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
		.SB_T0_NORTH_SB_IN_B16(Tile_X01_Y00_io2f_16),
		.SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B16),
		.SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B16),
		.SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B16),
		.SB_T0_WEST_SB_IN_B1(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_WEST_SB_IN_B16(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B16),
		.SB_T0_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B16(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B16),
		// .SB_T1_EAST_SB_IN_B1(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B1),
		// .SB_T1_EAST_SB_IN_B16(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B16),
		.SB_T1_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B16(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B16),
		.SB_T1_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
		.SB_T1_NORTH_SB_IN_B16(Tile_X01_Y00_io2f_16),
		.SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B16),
		.SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B16),
		.SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B16),
		.SB_T1_WEST_SB_IN_B1(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_WEST_SB_IN_B16(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B16),
		.SB_T1_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B16(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B16),
		// .SB_T2_EAST_SB_IN_B1(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B1),
		// .SB_T2_EAST_SB_IN_B16(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B16),
		.SB_T2_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B16(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B16),
		.SB_T2_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
		.SB_T2_NORTH_SB_IN_B16(Tile_X01_Y00_io2f_16),
		.SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B16),
		.SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B16),
		.SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B16),
		.SB_T2_WEST_SB_IN_B1(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_WEST_SB_IN_B16(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B16),
		.SB_T2_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B16(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B16),
		.clk(clk),
		.clk_out(Tile_X01_Y01_clk_out),
		.clk_pass_through(clk),
		.clk_pass_through_out_bot(Tile_X01_Y01_clk_pass_through_out_bot),
		.config_config_addr(config_1_config_addr),
		.config_config_data(config_1_config_data),
		.config_out_config_addr(Tile_X01_Y01_config_out_config_addr),
		.config_out_config_data(Tile_X01_Y01_config_out_config_data),
		.config_out_read(Tile_X01_Y01_config_out_read),
		.config_out_write(Tile_X01_Y01_config_out_write),
		.config_read(config_1_read),
		.config_write(config_1_write),
		.hi(Tile_X01_Y01_hi),
		.lo(Tile_X01_Y01_lo_unq1),
		.read_config_data(Tile_X01_Y01_read_config_data),
		.read_config_data_in(const_0_32_out),
		.reset(reset),
		.reset_out(Tile_X01_Y01_reset_out),
		.stall(stall[1]),
		.stall_out(Tile_X01_Y01_stall_out),
		.tile_id(Tile_X01_Y01_tile_id_in)
	);
	mantle_wire__typeBit8 Tile_X01_Y01_lo(
		.in(Tile_X01_Y01_lo_unq1),
		.out(Tile_X01_Y01_lo_out)
	);
	wire [15:0] Tile_X01_Y01_tile_id_out;
	assign Tile_X01_Y01_tile_id_out = {Tile_X01_Y01_lo_out[7], Tile_X01_Y01_lo_out[7:6], Tile_X01_Y01_lo_out[6:5], Tile_X01_Y01_lo_out[5:4], Tile_X01_Y01_hi[4], Tile_X01_Y01_lo_out[3], Tile_X01_Y01_lo_out[3:2], Tile_X01_Y01_lo_out[2:1], Tile_X01_Y01_lo_out[1:0], Tile_X01_Y01_hi[0]};
	mantle_wire__typeBitIn16 Tile_X01_Y01_tile_id(
		.in(Tile_X01_Y01_tile_id_in),
		.out(Tile_X01_Y01_tile_id_out)
	);
	Tile_PE Tile_X01_Y02(
		// .SB_T0_EAST_SB_IN_B1(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B1),
		// .SB_T0_EAST_SB_IN_B16(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B16),
		.SB_T0_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_EAST_SB_OUT_B16(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B16),
		.SB_T0_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_IN_B16(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B16),
		.SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B1),
		.SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B16),
		// .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B1),
		// .SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B16),
		.SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B1),
		.SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B16),
		.SB_T0_WEST_SB_IN_B1(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B1),
		.SB_T0_WEST_SB_IN_B16(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B16),
		.SB_T0_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B1),
		.SB_T0_WEST_SB_OUT_B16(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B16),
		// .SB_T1_EAST_SB_IN_B1(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B1),
		// .SB_T1_EAST_SB_IN_B16(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B16),
		.SB_T1_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_EAST_SB_OUT_B16(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B16),
		.SB_T1_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_IN_B16(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B16),
		.SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B1),
		.SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B16),
		// .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B1),
		// .SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B16),
		.SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B1),
		.SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B16),
		.SB_T1_WEST_SB_IN_B1(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B1),
		.SB_T1_WEST_SB_IN_B16(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B16),
		.SB_T1_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B1),
		.SB_T1_WEST_SB_OUT_B16(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B16),
		// .SB_T2_EAST_SB_IN_B1(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B1),
		// .SB_T2_EAST_SB_IN_B16(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B16),
		.SB_T2_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_EAST_SB_OUT_B16(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B16),
		.SB_T2_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_IN_B16(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B16),
		.SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B1),
		.SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B16),
		// .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B1),
		// .SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B16),
		.SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B1),
		.SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B16),
		.SB_T2_WEST_SB_IN_B1(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B1),
		.SB_T2_WEST_SB_IN_B16(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B16),
		.SB_T2_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B1),
		.SB_T2_WEST_SB_OUT_B16(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B16),
		.clk(Tile_X01_Y01_clk_out),
		.clk_out(Tile_X01_Y02_clk_out),
		.clk_pass_through(Tile_X01_Y01_clk_pass_through_out_bot),
		.clk_pass_through_out_bot(Tile_X01_Y02_clk_pass_through_out_bot),
		.config_config_addr(Tile_X01_Y01_config_out_config_addr),
		.config_config_data(Tile_X01_Y01_config_out_config_data),
		.config_out_config_addr(Tile_X01_Y02_config_out_config_addr),
		.config_out_config_data(Tile_X01_Y02_config_out_config_data),
		.config_out_read(Tile_X01_Y02_config_out_read),
		.config_out_write(Tile_X01_Y02_config_out_write),
		.config_read(Tile_X01_Y01_config_out_read),
		.config_write(Tile_X01_Y01_config_out_write),
		.hi(Tile_X01_Y02_hi),
		.lo(Tile_X01_Y02_lo_unq1),
		.read_config_data(Tile_X01_Y02_read_config_data),
		.read_config_data_in(Tile_X01_Y01_read_config_data),
		.reset(Tile_X01_Y01_reset_out),
		.reset_out(Tile_X01_Y02_reset_out),
		.stall(Tile_X01_Y01_stall_out),
		.stall_out(Tile_X01_Y02_stall_out),
		.tile_id(Tile_X01_Y02_tile_id_in)
	);
	mantle_wire__typeBit8 Tile_X01_Y02_lo(
		.in(Tile_X01_Y02_lo_unq1),
		.out(Tile_X01_Y02_lo_out)
	);
	wire [15:0] Tile_X01_Y02_tile_id_out;
	assign Tile_X01_Y02_tile_id_out = {Tile_X01_Y02_lo_out[7], Tile_X01_Y02_lo_out[7:6], Tile_X01_Y02_lo_out[6:5], Tile_X01_Y02_lo_out[5:4], Tile_X01_Y02_hi[4], Tile_X01_Y02_lo_out[3], Tile_X01_Y02_lo_out[3:2], Tile_X01_Y02_lo_out[2:1], Tile_X01_Y02_lo_out[1], Tile_X01_Y02_hi[1], Tile_X01_Y02_lo_out[0]};
	mantle_wire__typeBitIn16 Tile_X01_Y02_tile_id(
		.in(Tile_X01_Y02_tile_id_in),
		.out(Tile_X01_Y02_tile_id_out)
	);
	// Tile_PE Tile_X01_Y03(
	// 	.SB_T0_EAST_SB_IN_B1(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_IN_B16(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_IN_B16(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_IN_B16(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_IN_B16(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_IN_B16(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_IN_B16(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X01_Y02_clk_out),
	// 	.clk_out(Tile_X01_Y03_clk_out),
	// 	.clk_pass_through(Tile_X01_Y02_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X01_Y03_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X01_Y02_config_out_config_addr),
	// 	.config_config_data(Tile_X01_Y02_config_out_config_data),
	// 	.config_out_config_addr(Tile_X01_Y03_config_out_config_addr),
	// 	.config_out_config_data(Tile_X01_Y03_config_out_config_data),
	// 	.config_out_read(Tile_X01_Y03_config_out_read),
	// 	.config_out_write(Tile_X01_Y03_config_out_write),
	// 	.config_read(Tile_X01_Y02_config_out_read),
	// 	.config_write(Tile_X01_Y02_config_out_write),
	// 	.hi(Tile_X01_Y03_hi_unq1),
	// 	.lo(Tile_X01_Y03_lo_unq1),
	// 	.read_config_data(Tile_X01_Y03_read_config_data),
	// 	.read_config_data_in(Tile_X01_Y02_read_config_data),
	// 	.reset(Tile_X01_Y02_reset_out),
	// 	.reset_out(Tile_X01_Y03_reset_out),
	// 	.stall(Tile_X01_Y02_stall_out),
	// 	.stall_out(Tile_X01_Y03_stall_out),
	// 	.tile_id(Tile_X01_Y03_tile_id_in)
	// );
	// mantle_wire__typeBit9 Tile_X01_Y03_hi(
	// 	.in(Tile_X01_Y03_hi_unq1),
	// 	.out(Tile_X01_Y03_hi_out)
	// );
	// mantle_wire__typeBit8 Tile_X01_Y03_lo(
	// 	.in(Tile_X01_Y03_lo_unq1),
	// 	.out(Tile_X01_Y03_lo_out)
	// );
	// wire [15:0] Tile_X01_Y03_tile_id_out;
	// assign Tile_X01_Y03_tile_id_out = {Tile_X01_Y03_lo_out[7], Tile_X01_Y03_lo_out[7:6], Tile_X01_Y03_lo_out[6:5], Tile_X01_Y03_lo_out[5:4], Tile_X01_Y03_hi_out[4], Tile_X01_Y03_lo_out[3], Tile_X01_Y03_lo_out[3:2], Tile_X01_Y03_lo_out[2:1], Tile_X01_Y03_lo_out[1], Tile_X01_Y03_hi_out[1:0]};
	// mantle_wire__typeBitIn16 Tile_X01_Y03_tile_id(
	// 	.in(Tile_X01_Y03_tile_id_in),
	// 	.out(Tile_X01_Y03_tile_id_out)
	// );
	// Tile_PE Tile_X01_Y04(
	// 	.SB_T0_EAST_SB_IN_B1(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_IN_B16(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y05_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y05_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_IN_B16(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_IN_B16(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y05_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y05_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_IN_B16(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_IN_B16(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y05_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y05_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_IN_B16(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X01_Y03_clk_out),
	// 	.clk_out(Tile_X01_Y04_clk_out),
	// 	.clk_pass_through(Tile_X01_Y03_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X01_Y04_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X01_Y03_config_out_config_addr),
	// 	.config_config_data(Tile_X01_Y03_config_out_config_data),
	// 	.config_out_config_addr(Tile_X01_Y04_config_out_config_addr),
	// 	.config_out_config_data(Tile_X01_Y04_config_out_config_data),
	// 	.config_out_read(Tile_X01_Y04_config_out_read),
	// 	.config_out_write(Tile_X01_Y04_config_out_write),
	// 	.config_read(Tile_X01_Y03_config_out_read),
	// 	.config_write(Tile_X01_Y03_config_out_write),
	// 	.hi(Tile_X01_Y04_hi),
	// 	.lo(Tile_X01_Y04_lo_unq1),
	// 	.read_config_data(Tile_X01_Y04_read_config_data),
	// 	.read_config_data_in(Tile_X01_Y03_read_config_data),
	// 	.reset(Tile_X01_Y03_reset_out),
	// 	.reset_out(Tile_X01_Y04_reset_out),
	// 	.stall(Tile_X01_Y03_stall_out),
	// 	.stall_out(Tile_X01_Y04_stall_out),
	// 	.tile_id(Tile_X01_Y04_tile_id_in)
	// );
	// mantle_wire__typeBit8 Tile_X01_Y04_lo(
	// 	.in(Tile_X01_Y04_lo_unq1),
	// 	.out(Tile_X01_Y04_lo_out)
	// );
	// wire [15:0] Tile_X01_Y04_tile_id_out;
	// assign Tile_X01_Y04_tile_id_out = {Tile_X01_Y04_lo_out[7], Tile_X01_Y04_lo_out[7:6], Tile_X01_Y04_lo_out[6:5], Tile_X01_Y04_lo_out[5:4], Tile_X01_Y04_hi[4], Tile_X01_Y04_lo_out[3], Tile_X01_Y04_lo_out[3:2], Tile_X01_Y04_lo_out[2:1], Tile_X01_Y04_hi[1], Tile_X01_Y04_lo_out[0], Tile_X01_Y04_lo_out[0]};
	// mantle_wire__typeBitIn16 Tile_X01_Y04_tile_id(
	// 	.in(Tile_X01_Y04_tile_id_in),
	// 	.out(Tile_X01_Y04_tile_id_out)
	// );
	// Tile_MemCore Tile_X01_Y05(
	// 	.SB_T0_EAST_SB_IN_B1(Tile_X02_Y05_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_IN_B16(Tile_X02_Y05_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X01_Y05_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X01_Y05_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y05_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y05_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y06_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y06_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y05_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y05_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(Tile_X00_Y05_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_IN_B16(Tile_X00_Y05_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X01_Y05_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X01_Y05_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(Tile_X02_Y05_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_IN_B16(Tile_X02_Y05_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X01_Y05_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X01_Y05_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y05_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y05_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y06_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y06_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y05_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y05_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(Tile_X00_Y05_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_IN_B16(Tile_X00_Y05_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X01_Y05_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X01_Y05_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(Tile_X02_Y05_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_IN_B16(Tile_X02_Y05_SB_T2_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X01_Y05_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X01_Y05_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y05_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y05_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y06_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y06_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y05_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y05_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(Tile_X00_Y05_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_IN_B16(Tile_X00_Y05_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X01_Y05_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X01_Y05_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X01_Y04_clk_out),
	// 	.clk_out(Tile_X01_Y05_clk_out),
	// 	.clk_pass_through(Tile_X01_Y04_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X01_Y05_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X01_Y04_config_out_config_addr),
	// 	.config_config_data(Tile_X01_Y04_config_out_config_data),
	// 	.config_out_config_addr(Tile_X01_Y05_config_out_config_addr),
	// 	.config_out_config_data(Tile_X01_Y05_config_out_config_data),
	// 	.config_out_read(Tile_X01_Y05_config_out_read),
	// 	.config_out_write(Tile_X01_Y05_config_out_write),
	// 	.config_read(Tile_X01_Y04_config_out_read),
	// 	.config_write(Tile_X01_Y04_config_out_write),
	// 	.hi(Tile_X01_Y05_hi),
	// 	.lo(Tile_X01_Y05_lo_unq1),
	// 	.read_config_data(Tile_X01_Y05_read_config_data),
	// 	.read_config_data_in(Tile_X01_Y04_read_config_data),
	// 	.reset(Tile_X01_Y04_reset_out),
	// 	.reset_out(Tile_X01_Y05_reset_out),
	// 	.stall(Tile_X01_Y04_stall_out),
	// 	.stall_out(Tile_X01_Y05_stall_out),
	// 	.tile_id(Tile_X01_Y05_tile_id_in)
	// );
	// mantle_wire__typeBit8 Tile_X01_Y05_lo(
	// 	.in(Tile_X01_Y05_lo_unq1),
	// 	.out(Tile_X01_Y05_lo_out)
	// );
	// wire [15:0] Tile_X01_Y05_tile_id_out;
	// assign Tile_X01_Y05_tile_id_out = {Tile_X01_Y05_lo_out[7], Tile_X01_Y05_lo_out[7:6], Tile_X01_Y05_lo_out[6:5], Tile_X01_Y05_lo_out[5:4], Tile_X01_Y05_hi[4], Tile_X01_Y05_lo_out[3], Tile_X01_Y05_lo_out[3:2], Tile_X01_Y05_lo_out[2:1], Tile_X01_Y05_hi[1], Tile_X01_Y05_lo_out[0], Tile_X01_Y05_hi[0]};
	// mantle_wire__typeBitIn16 Tile_X01_Y05_tile_id(
	// 	.in(Tile_X01_Y05_tile_id_in),
	// 	.out(Tile_X01_Y05_tile_id_out)
	// );
	// Tile_PE Tile_X01_Y06(
	// 	.SB_T0_EAST_SB_IN_B1(Tile_X02_Y06_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_IN_B16(Tile_X02_Y06_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X01_Y06_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X01_Y06_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X01_Y05_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X01_Y05_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y06_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y06_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y07_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y07_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y06_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y06_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(Tile_X00_Y06_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_IN_B16(Tile_X00_Y06_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X01_Y06_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X01_Y06_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(Tile_X02_Y06_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_IN_B16(Tile_X02_Y06_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X01_Y06_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X01_Y06_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X01_Y05_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X01_Y05_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y06_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y06_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y07_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y07_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y06_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y06_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(Tile_X00_Y06_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_IN_B16(Tile_X00_Y06_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X01_Y06_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X01_Y06_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(Tile_X02_Y06_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_IN_B16(Tile_X02_Y06_SB_T2_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X01_Y06_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X01_Y06_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X01_Y05_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X01_Y05_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y06_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y06_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y07_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y07_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y06_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y06_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(Tile_X00_Y06_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_IN_B16(Tile_X00_Y06_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X01_Y06_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X01_Y06_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X01_Y05_clk_out),
	// 	.clk_out(Tile_X01_Y06_clk_out),
	// 	.clk_pass_through(Tile_X01_Y05_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X01_Y06_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X01_Y05_config_out_config_addr),
	// 	.config_config_data(Tile_X01_Y05_config_out_config_data),
	// 	.config_out_config_addr(Tile_X01_Y06_config_out_config_addr),
	// 	.config_out_config_data(Tile_X01_Y06_config_out_config_data),
	// 	.config_out_read(Tile_X01_Y06_config_out_read),
	// 	.config_out_write(Tile_X01_Y06_config_out_write),
	// 	.config_read(Tile_X01_Y05_config_out_read),
	// 	.config_write(Tile_X01_Y05_config_out_write),
	// 	.hi(Tile_X01_Y06_hi),
	// 	.lo(Tile_X01_Y06_lo_unq1),
	// 	.read_config_data(Tile_X01_Y06_read_config_data),
	// 	.read_config_data_in(Tile_X01_Y05_read_config_data),
	// 	.reset(Tile_X01_Y05_reset_out),
	// 	.reset_out(Tile_X01_Y06_reset_out),
	// 	.stall(Tile_X01_Y05_stall_out),
	// 	.stall_out(Tile_X01_Y06_stall_out),
	// 	.tile_id(Tile_X01_Y06_tile_id_in)
	// );
	// mantle_wire__typeBit8 Tile_X01_Y06_lo(
	// 	.in(Tile_X01_Y06_lo_unq1),
	// 	.out(Tile_X01_Y06_lo_out)
	// );
	// wire [15:0] Tile_X01_Y06_tile_id_out;
	// assign Tile_X01_Y06_tile_id_out = {Tile_X01_Y06_lo_out[7], Tile_X01_Y06_lo_out[7:6], Tile_X01_Y06_lo_out[6:5], Tile_X01_Y06_lo_out[5:4], Tile_X01_Y06_hi[4], Tile_X01_Y06_lo_out[3], Tile_X01_Y06_lo_out[3:2], Tile_X01_Y06_lo_out[2:1], Tile_X01_Y06_hi[1], Tile_X01_Y06_hi[1], Tile_X01_Y06_lo_out[0]};
	// mantle_wire__typeBitIn16 Tile_X01_Y06_tile_id(
	// 	.in(Tile_X01_Y06_tile_id_in),
	// 	.out(Tile_X01_Y06_tile_id_out)
	// );
	// Tile_PE Tile_X01_Y07(
	// 	.SB_T0_EAST_SB_IN_B1(Tile_X02_Y07_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_IN_B16(Tile_X02_Y07_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X01_Y07_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X01_Y07_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X01_Y06_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X01_Y06_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y07_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y07_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y08_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y08_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y07_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y07_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(Tile_X00_Y07_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_IN_B16(Tile_X00_Y07_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X01_Y07_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X01_Y07_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(Tile_X02_Y07_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_IN_B16(Tile_X02_Y07_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X01_Y07_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X01_Y07_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X01_Y06_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X01_Y06_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y07_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y07_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y08_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y08_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y07_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y07_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(Tile_X00_Y07_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_IN_B16(Tile_X00_Y07_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X01_Y07_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X01_Y07_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(Tile_X02_Y07_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_IN_B16(Tile_X02_Y07_SB_T2_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X01_Y07_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X01_Y07_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X01_Y06_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X01_Y06_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y07_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y07_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y08_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y08_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y07_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y07_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(Tile_X00_Y07_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_IN_B16(Tile_X00_Y07_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X01_Y07_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X01_Y07_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X01_Y06_clk_out),
	// 	.clk_out(Tile_X01_Y07_clk_out),
	// 	.clk_pass_through(Tile_X01_Y06_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X01_Y07_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X01_Y06_config_out_config_addr),
	// 	.config_config_data(Tile_X01_Y06_config_out_config_data),
	// 	.config_out_config_addr(Tile_X01_Y07_config_out_config_addr),
	// 	.config_out_config_data(Tile_X01_Y07_config_out_config_data),
	// 	.config_out_read(Tile_X01_Y07_config_out_read),
	// 	.config_out_write(Tile_X01_Y07_config_out_write),
	// 	.config_read(Tile_X01_Y06_config_out_read),
	// 	.config_write(Tile_X01_Y06_config_out_write),
	// 	.hi(Tile_X01_Y07_hi_unq1),
	// 	.lo(Tile_X01_Y07_lo_unq1),
	// 	.read_config_data(Tile_X01_Y07_read_config_data),
	// 	.read_config_data_in(Tile_X01_Y06_read_config_data),
	// 	.reset(Tile_X01_Y06_reset_out),
	// 	.reset_out(Tile_X01_Y07_reset_out),
	// 	.stall(Tile_X01_Y06_stall_out),
	// 	.stall_out(Tile_X01_Y07_stall_out),
	// 	.tile_id(Tile_X01_Y07_tile_id_in)
	// );
	// mantle_wire__typeBit9 Tile_X01_Y07_hi(
	// 	.in(Tile_X01_Y07_hi_unq1),
	// 	.out(Tile_X01_Y07_hi_out)
	// );
	// mantle_wire__typeBit8 Tile_X01_Y07_lo(
	// 	.in(Tile_X01_Y07_lo_unq1),
	// 	.out(Tile_X01_Y07_lo_out)
	// );
	// wire [15:0] Tile_X01_Y07_tile_id_out;
	// assign Tile_X01_Y07_tile_id_out = {Tile_X01_Y07_lo_out[7], Tile_X01_Y07_lo_out[7:6], Tile_X01_Y07_lo_out[6:5], Tile_X01_Y07_lo_out[5:4], Tile_X01_Y07_hi_out[4], Tile_X01_Y07_lo_out[3], Tile_X01_Y07_lo_out[3:2], Tile_X01_Y07_lo_out[2:1], Tile_X01_Y07_hi_out[1], Tile_X01_Y07_hi_out[1:0]};
	// mantle_wire__typeBitIn16 Tile_X01_Y07_tile_id(
	// 	.in(Tile_X01_Y07_tile_id_in),
	// 	.out(Tile_X01_Y07_tile_id_out)
	// );
	// Tile_PE Tile_X01_Y08(
	// 	.SB_T0_EAST_SB_IN_B1(Tile_X02_Y08_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_IN_B16(Tile_X02_Y08_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X01_Y08_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X01_Y08_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X01_Y07_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X01_Y07_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y08_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y08_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
	// 	.SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y08_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y08_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(Tile_X00_Y08_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_IN_B16(Tile_X00_Y08_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X01_Y08_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X01_Y08_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(Tile_X02_Y08_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_IN_B16(Tile_X02_Y08_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X01_Y08_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X01_Y08_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X01_Y07_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X01_Y07_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y08_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y08_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
	// 	.SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y08_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y08_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(Tile_X00_Y08_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_IN_B16(Tile_X00_Y08_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X01_Y08_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X01_Y08_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(Tile_X02_Y08_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_IN_B16(Tile_X02_Y08_SB_T2_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X01_Y08_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X01_Y08_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X01_Y07_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X01_Y07_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y08_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y08_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
	// 	.SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y08_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y08_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(Tile_X00_Y08_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_IN_B16(Tile_X00_Y08_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X01_Y08_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X01_Y08_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X01_Y07_clk_out),
	// 	.clk_out(Tile_X01_Y08_clk_out),
	// 	.clk_pass_through(Tile_X01_Y07_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X01_Y08_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X01_Y07_config_out_config_addr),
	// 	.config_config_data(Tile_X01_Y07_config_out_config_data),
	// 	.config_out_config_addr(Tile_X01_Y08_config_out_config_addr),
	// 	.config_out_config_data(Tile_X01_Y08_config_out_config_data),
	// 	.config_out_read(Tile_X01_Y08_config_out_read),
	// 	.config_out_write(Tile_X01_Y08_config_out_write),
	// 	.config_read(Tile_X01_Y07_config_out_read),
	// 	.config_write(Tile_X01_Y07_config_out_write),
	// 	.hi(Tile_X01_Y08_hi),
	// 	.lo(Tile_X01_Y08_lo_unq1),
	// 	.read_config_data(Tile_X01_Y08_read_config_data),
	// 	.read_config_data_in(Tile_X01_Y07_read_config_data),
	// 	.reset(Tile_X01_Y07_reset_out),
	// 	.reset_out(Tile_X01_Y08_reset_out),
	// 	.stall(Tile_X01_Y07_stall_out),
	// 	.stall_out(Tile_X01_Y08_stall_out),
	// 	.tile_id(Tile_X01_Y08_tile_id_in)
	// );
	// mantle_wire__typeBit8 Tile_X01_Y08_lo(
	// 	.in(Tile_X01_Y08_lo_unq1),
	// 	.out(Tile_X01_Y08_lo_out)
	// );
	// wire [15:0] Tile_X01_Y08_tile_id_out;
	// assign Tile_X01_Y08_tile_id_out = {Tile_X01_Y08_lo_out[7], Tile_X01_Y08_lo_out[7:6], Tile_X01_Y08_lo_out[6:5], Tile_X01_Y08_lo_out[5:4], Tile_X01_Y08_hi[4], Tile_X01_Y08_lo_out[3], Tile_X01_Y08_lo_out[3:2], Tile_X01_Y08_lo_out[2], Tile_X01_Y08_hi[2], Tile_X01_Y08_lo_out[1:0], Tile_X01_Y08_lo_out[0]};
	// mantle_wire__typeBitIn16 Tile_X01_Y08_tile_id(
	// 	.in(Tile_X01_Y08_tile_id_in),
	// 	.out(Tile_X01_Y08_tile_id_out)
	// );
	// wire [15:0] Tile_X02_Y00_tile_id;
	// assign Tile_X02_Y00_tile_id = {Tile_X02_Y00_lo[7], Tile_X02_Y00_lo[7:6], Tile_X02_Y00_lo[6:5], Tile_X02_Y00_lo[5], Tile_X02_Y00_hi[5], Tile_X02_Y00_lo[4:3], Tile_X02_Y00_lo[3:2], Tile_X02_Y00_lo[2:1], Tile_X02_Y00_lo[1:0], Tile_X02_Y00_lo[0]};
	// Tile_io_core Tile_X02_Y00(
	// 	.tile_id(Tile_X02_Y00_tile_id),
	// 	.glb2io_1(glb2io_1_X02_Y00),
	// 	.f2io_1(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B1),
	// 	.io2glb_1(Tile_X02_Y00_io2glb_1),
	// 	.io2f_1(Tile_X02_Y00_io2f_1),
	// 	.glb2io_16(glb2io_16_X02_Y00),
	// 	.f2io_16(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B16),
	// 	.io2glb_16(Tile_X02_Y00_io2glb_16),
	// 	.io2f_16(Tile_X02_Y00_io2f_16),
	// 	.hi(Tile_X02_Y00_hi),
	// 	.lo(Tile_X02_Y00_lo)
	// );
	// Tile_MemCore Tile_X02_Y01(
	// 	.SB_T0_EAST_SB_IN_B1(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_IN_B16(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X02_Y00_io2f_16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B16),
	// 	// .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B1),
	// 	// .SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B16),
	// 	// .SB_T0_WEST_SB_IN_B1(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B1),
	// 	// .SB_T0_WEST_SB_IN_B16(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_IN_B16(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X02_Y00_io2f_16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B16),
	// 	// .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B1),
	// 	// .SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B16),
	// 	// .SB_T1_WEST_SB_IN_B1(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B1),
	// 	// .SB_T1_WEST_SB_IN_B16(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_IN_B16(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X02_Y00_io2f_16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B16),
	// 	// .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B1),
	// 	// .SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B16),
	// 	// .SB_T2_WEST_SB_IN_B1(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B1),
	// 	// .SB_T2_WEST_SB_IN_B16(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(clk),
	// 	.clk_out(Tile_X02_Y01_clk_out),
	// 	.clk_pass_through(clk),
	// 	.clk_pass_through_out_bot(Tile_X02_Y01_clk_pass_through_out_bot),
	// 	.config_config_addr(config_2_config_addr),
	// 	.config_config_data(config_2_config_data),
	// 	.config_out_config_addr(Tile_X02_Y01_config_out_config_addr),
	// 	.config_out_config_data(Tile_X02_Y01_config_out_config_data),
	// 	.config_out_read(Tile_X02_Y01_config_out_read),
	// 	.config_out_write(Tile_X02_Y01_config_out_write),
	// 	.config_read(config_2_read),
	// 	.config_write(config_2_write),
	// 	.hi(Tile_X02_Y01_hi),
	// 	.lo(Tile_X02_Y01_lo_unq1),
	// 	.read_config_data(Tile_X02_Y01_read_config_data),
	// 	.read_config_data_in(const_0_32_out),
	// 	.reset(reset),
	// 	.reset_out(Tile_X02_Y01_reset_out),
	// 	.stall(stall[2]),
	// 	.stall_out(Tile_X02_Y01_stall_out),
	// 	.tile_id(Tile_X02_Y01_tile_id_in)
	// );
	// mantle_wire__typeBit8 Tile_X02_Y01_lo(
	// 	.in(Tile_X02_Y01_lo_unq1),
	// 	.out(Tile_X02_Y01_lo_out)
	// );
	// wire [15:0] Tile_X02_Y01_tile_id_out;
	// assign Tile_X02_Y01_tile_id_out = {Tile_X02_Y01_lo_out[7], Tile_X02_Y01_lo_out[7:6], Tile_X02_Y01_lo_out[6:5], Tile_X02_Y01_lo_out[5], Tile_X02_Y01_hi[5], Tile_X02_Y01_lo_out[4:3], Tile_X02_Y01_lo_out[3:2], Tile_X02_Y01_lo_out[2:1], Tile_X02_Y01_lo_out[1:0], Tile_X02_Y01_hi[0]};
	// mantle_wire__typeBitIn16 Tile_X02_Y01_tile_id(
	// 	.in(Tile_X02_Y01_tile_id_in),
	// 	.out(Tile_X02_Y01_tile_id_out)
	// );
	// Tile_PE Tile_X02_Y02(
	// 	.SB_T0_EAST_SB_IN_B1(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_IN_B16(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B16),
	// 	// .SB_T0_WEST_SB_IN_B1(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B1),
	// 	// .SB_T0_WEST_SB_IN_B16(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_IN_B16(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B16),
	// 	// .SB_T1_WEST_SB_IN_B1(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B1),
	// 	// .SB_T1_WEST_SB_IN_B16(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_IN_B16(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B16),
	// 	// .SB_T2_WEST_SB_IN_B1(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B1),
	// 	// .SB_T2_WEST_SB_IN_B16(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X02_Y01_clk_out),
	// 	.clk_out(Tile_X02_Y02_clk_out),
	// 	.clk_pass_through(Tile_X02_Y01_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X02_Y02_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X02_Y01_config_out_config_addr),
	// 	.config_config_data(Tile_X02_Y01_config_out_config_data),
	// 	.config_out_config_addr(Tile_X02_Y02_config_out_config_addr),
	// 	.config_out_config_data(Tile_X02_Y02_config_out_config_data),
	// 	.config_out_read(Tile_X02_Y02_config_out_read),
	// 	.config_out_write(Tile_X02_Y02_config_out_write),
	// 	.config_read(Tile_X02_Y01_config_out_read),
	// 	.config_write(Tile_X02_Y01_config_out_write),
	// 	.hi(Tile_X02_Y02_hi),
	// 	.lo(Tile_X02_Y02_lo_unq1),
	// 	.read_config_data(Tile_X02_Y02_read_config_data),
	// 	.read_config_data_in(Tile_X02_Y01_read_config_data),
	// 	.reset(Tile_X02_Y01_reset_out),
	// 	.reset_out(Tile_X02_Y02_reset_out),
	// 	.stall(Tile_X02_Y01_stall_out),
	// 	.stall_out(Tile_X02_Y02_stall_out),
	// 	.tile_id(Tile_X02_Y02_tile_id_in)
	// );
	// mantle_wire__typeBit8 Tile_X02_Y02_lo(
	// 	.in(Tile_X02_Y02_lo_unq1),
	// 	.out(Tile_X02_Y02_lo_out)
	// );
	// wire [15:0] Tile_X02_Y02_tile_id_out;
	// assign Tile_X02_Y02_tile_id_out = {Tile_X02_Y02_lo_out[7], Tile_X02_Y02_lo_out[7:6], Tile_X02_Y02_lo_out[6:5], Tile_X02_Y02_lo_out[5], Tile_X02_Y02_hi[5], Tile_X02_Y02_lo_out[4:3], Tile_X02_Y02_lo_out[3:2], Tile_X02_Y02_lo_out[2:1], Tile_X02_Y02_lo_out[1], Tile_X02_Y02_hi[1], Tile_X02_Y02_lo_out[0]};
	// mantle_wire__typeBitIn16 Tile_X02_Y02_tile_id(
	// 	.in(Tile_X02_Y02_tile_id_in),
	// 	.out(Tile_X02_Y02_tile_id_out)
	// );
	// Tile_PE Tile_X02_Y03(
	// 	.SB_T0_EAST_SB_IN_B1(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_IN_B16(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_IN_B16(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_IN_B16(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_IN_B16(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_IN_B16(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_IN_B16(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X02_Y02_clk_out),
	// 	.clk_out(Tile_X02_Y03_clk_out),
	// 	.clk_pass_through(Tile_X02_Y02_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X02_Y03_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X02_Y02_config_out_config_addr),
	// 	.config_config_data(Tile_X02_Y02_config_out_config_data),
	// 	.config_out_config_addr(Tile_X02_Y03_config_out_config_addr),
	// 	.config_out_config_data(Tile_X02_Y03_config_out_config_data),
	// 	.config_out_read(Tile_X02_Y03_config_out_read),
	// 	.config_out_write(Tile_X02_Y03_config_out_write),
	// 	.config_read(Tile_X02_Y02_config_out_read),
	// 	.config_write(Tile_X02_Y02_config_out_write),
	// 	.hi(Tile_X02_Y03_hi_unq1),
	// 	.lo(Tile_X02_Y03_lo_unq1),
	// 	.read_config_data(Tile_X02_Y03_read_config_data),
	// 	.read_config_data_in(Tile_X02_Y02_read_config_data),
	// 	.reset(Tile_X02_Y02_reset_out),
	// 	.reset_out(Tile_X02_Y03_reset_out),
	// 	.stall(Tile_X02_Y02_stall_out),
	// 	.stall_out(Tile_X02_Y03_stall_out),
	// 	.tile_id(Tile_X02_Y03_tile_id_in)
	// );
	// mantle_wire__typeBit9 Tile_X02_Y03_hi(
	// 	.in(Tile_X02_Y03_hi_unq1),
	// 	.out(Tile_X02_Y03_hi_out)
	// );
	// mantle_wire__typeBit8 Tile_X02_Y03_lo(
	// 	.in(Tile_X02_Y03_lo_unq1),
	// 	.out(Tile_X02_Y03_lo_out)
	// );
	// wire [15:0] Tile_X02_Y03_tile_id_out;
	// assign Tile_X02_Y03_tile_id_out = {Tile_X02_Y03_lo_out[7], Tile_X02_Y03_lo_out[7:6], Tile_X02_Y03_lo_out[6:5], Tile_X02_Y03_lo_out[5], Tile_X02_Y03_hi_out[5], Tile_X02_Y03_lo_out[4:3], Tile_X02_Y03_lo_out[3:2], Tile_X02_Y03_lo_out[2:1], Tile_X02_Y03_lo_out[1], Tile_X02_Y03_hi_out[1:0]};
	// mantle_wire__typeBitIn16 Tile_X02_Y03_tile_id(
	// 	.in(Tile_X02_Y03_tile_id_in),
	// 	.out(Tile_X02_Y03_tile_id_out)
	// );
	// Tile_PE Tile_X02_Y04(
	// 	.SB_T0_EAST_SB_IN_B1(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_IN_B16(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y05_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y05_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_IN_B16(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_IN_B16(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y05_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y05_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_IN_B16(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_IN_B16(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y05_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y05_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_IN_B16(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X02_Y03_clk_out),
	// 	.clk_out(Tile_X02_Y04_clk_out),
	// 	.clk_pass_through(Tile_X02_Y03_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X02_Y04_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X02_Y03_config_out_config_addr),
	// 	.config_config_data(Tile_X02_Y03_config_out_config_data),
	// 	.config_out_config_addr(Tile_X02_Y04_config_out_config_addr),
	// 	.config_out_config_data(Tile_X02_Y04_config_out_config_data),
	// 	.config_out_read(Tile_X02_Y04_config_out_read),
	// 	.config_out_write(Tile_X02_Y04_config_out_write),
	// 	.config_read(Tile_X02_Y03_config_out_read),
	// 	.config_write(Tile_X02_Y03_config_out_write),
	// 	.hi(Tile_X02_Y04_hi),
	// 	.lo(Tile_X02_Y04_lo_unq1),
	// 	.read_config_data(Tile_X02_Y04_read_config_data),
	// 	.read_config_data_in(Tile_X02_Y03_read_config_data),
	// 	.reset(Tile_X02_Y03_reset_out),
	// 	.reset_out(Tile_X02_Y04_reset_out),
	// 	.stall(Tile_X02_Y03_stall_out),
	// 	.stall_out(Tile_X02_Y04_stall_out),
	// 	.tile_id(Tile_X02_Y04_tile_id_in)
	// );
	// mantle_wire__typeBit8 Tile_X02_Y04_lo(
	// 	.in(Tile_X02_Y04_lo_unq1),
	// 	.out(Tile_X02_Y04_lo_out)
	// );
	// wire [15:0] Tile_X02_Y04_tile_id_out;
	// assign Tile_X02_Y04_tile_id_out = {Tile_X02_Y04_lo_out[7], Tile_X02_Y04_lo_out[7:6], Tile_X02_Y04_lo_out[6:5], Tile_X02_Y04_lo_out[5], Tile_X02_Y04_hi[5], Tile_X02_Y04_lo_out[4:3], Tile_X02_Y04_lo_out[3:2], Tile_X02_Y04_lo_out[2:1], Tile_X02_Y04_hi[1], Tile_X02_Y04_lo_out[0], Tile_X02_Y04_lo_out[0]};
	// mantle_wire__typeBitIn16 Tile_X02_Y04_tile_id(
	// 	.in(Tile_X02_Y04_tile_id_in),
	// 	.out(Tile_X02_Y04_tile_id_out)
	// );
	// Tile_MemCore Tile_X02_Y05(
	// 	.SB_T0_EAST_SB_IN_B1(Tile_X03_Y05_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_IN_B16(Tile_X03_Y05_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X02_Y05_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X02_Y05_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y05_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y05_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y06_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y06_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y05_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y05_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(Tile_X01_Y05_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_IN_B16(Tile_X01_Y05_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X02_Y05_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X02_Y05_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(Tile_X03_Y05_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_IN_B16(Tile_X03_Y05_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X02_Y05_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X02_Y05_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y05_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y05_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y06_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y06_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y05_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y05_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(Tile_X01_Y05_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_IN_B16(Tile_X01_Y05_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X02_Y05_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X02_Y05_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(Tile_X03_Y05_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_IN_B16(Tile_X03_Y05_SB_T2_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X02_Y05_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X02_Y05_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y05_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y05_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y06_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y06_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y05_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y05_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(Tile_X01_Y05_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_IN_B16(Tile_X01_Y05_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X02_Y05_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X02_Y05_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X02_Y04_clk_out),
	// 	.clk_out(Tile_X02_Y05_clk_out),
	// 	.clk_pass_through(Tile_X02_Y04_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X02_Y05_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X02_Y04_config_out_config_addr),
	// 	.config_config_data(Tile_X02_Y04_config_out_config_data),
	// 	.config_out_config_addr(Tile_X02_Y05_config_out_config_addr),
	// 	.config_out_config_data(Tile_X02_Y05_config_out_config_data),
	// 	.config_out_read(Tile_X02_Y05_config_out_read),
	// 	.config_out_write(Tile_X02_Y05_config_out_write),
	// 	.config_read(Tile_X02_Y04_config_out_read),
	// 	.config_write(Tile_X02_Y04_config_out_write),
	// 	.hi(Tile_X02_Y05_hi),
	// 	.lo(Tile_X02_Y05_lo_unq1),
	// 	.read_config_data(Tile_X02_Y05_read_config_data),
	// 	.read_config_data_in(Tile_X02_Y04_read_config_data),
	// 	.reset(Tile_X02_Y04_reset_out),
	// 	.reset_out(Tile_X02_Y05_reset_out),
	// 	.stall(Tile_X02_Y04_stall_out),
	// 	.stall_out(Tile_X02_Y05_stall_out),
	// 	.tile_id(Tile_X02_Y05_tile_id_in)
	// );
	// mantle_wire__typeBit8 Tile_X02_Y05_lo(
	// 	.in(Tile_X02_Y05_lo_unq1),
	// 	.out(Tile_X02_Y05_lo_out)
	// );
	// wire [15:0] Tile_X02_Y05_tile_id_out;
	// assign Tile_X02_Y05_tile_id_out = {Tile_X02_Y05_lo_out[7], Tile_X02_Y05_lo_out[7:6], Tile_X02_Y05_lo_out[6:5], Tile_X02_Y05_lo_out[5], Tile_X02_Y05_hi[5], Tile_X02_Y05_lo_out[4:3], Tile_X02_Y05_lo_out[3:2], Tile_X02_Y05_lo_out[2:1], Tile_X02_Y05_hi[1], Tile_X02_Y05_lo_out[0], Tile_X02_Y05_hi[0]};
	// mantle_wire__typeBitIn16 Tile_X02_Y05_tile_id(
	// 	.in(Tile_X02_Y05_tile_id_in),
	// 	.out(Tile_X02_Y05_tile_id_out)
	// );
	// Tile_PE Tile_X02_Y06(
	// 	.SB_T0_EAST_SB_IN_B1(Tile_X03_Y06_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_IN_B16(Tile_X03_Y06_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X02_Y06_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X02_Y06_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X02_Y05_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X02_Y05_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y06_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y06_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y07_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y07_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y06_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y06_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(Tile_X01_Y06_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_IN_B16(Tile_X01_Y06_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X02_Y06_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X02_Y06_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(Tile_X03_Y06_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_IN_B16(Tile_X03_Y06_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X02_Y06_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X02_Y06_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X02_Y05_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X02_Y05_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y06_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y06_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y07_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y07_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y06_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y06_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(Tile_X01_Y06_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_IN_B16(Tile_X01_Y06_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X02_Y06_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X02_Y06_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(Tile_X03_Y06_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_IN_B16(Tile_X03_Y06_SB_T2_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X02_Y06_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X02_Y06_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X02_Y05_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X02_Y05_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y06_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y06_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y07_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y07_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y06_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y06_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(Tile_X01_Y06_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_IN_B16(Tile_X01_Y06_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X02_Y06_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X02_Y06_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X02_Y05_clk_out),
	// 	.clk_out(Tile_X02_Y06_clk_out),
	// 	.clk_pass_through(Tile_X02_Y05_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X02_Y06_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X02_Y05_config_out_config_addr),
	// 	.config_config_data(Tile_X02_Y05_config_out_config_data),
	// 	.config_out_config_addr(Tile_X02_Y06_config_out_config_addr),
	// 	.config_out_config_data(Tile_X02_Y06_config_out_config_data),
	// 	.config_out_read(Tile_X02_Y06_config_out_read),
	// 	.config_out_write(Tile_X02_Y06_config_out_write),
	// 	.config_read(Tile_X02_Y05_config_out_read),
	// 	.config_write(Tile_X02_Y05_config_out_write),
	// 	.hi(Tile_X02_Y06_hi),
	// 	.lo(Tile_X02_Y06_lo_unq1),
	// 	.read_config_data(Tile_X02_Y06_read_config_data),
	// 	.read_config_data_in(Tile_X02_Y05_read_config_data),
	// 	.reset(Tile_X02_Y05_reset_out),
	// 	.reset_out(Tile_X02_Y06_reset_out),
	// 	.stall(Tile_X02_Y05_stall_out),
	// 	.stall_out(Tile_X02_Y06_stall_out),
	// 	.tile_id(Tile_X02_Y06_tile_id_in)
	// );
	// mantle_wire__typeBit8 Tile_X02_Y06_lo(
	// 	.in(Tile_X02_Y06_lo_unq1),
	// 	.out(Tile_X02_Y06_lo_out)
	// );
	// wire [15:0] Tile_X02_Y06_tile_id_out;
	// assign Tile_X02_Y06_tile_id_out = {Tile_X02_Y06_lo_out[7], Tile_X02_Y06_lo_out[7:6], Tile_X02_Y06_lo_out[6:5], Tile_X02_Y06_lo_out[5], Tile_X02_Y06_hi[5], Tile_X02_Y06_lo_out[4:3], Tile_X02_Y06_lo_out[3:2], Tile_X02_Y06_lo_out[2:1], Tile_X02_Y06_hi[1], Tile_X02_Y06_hi[1], Tile_X02_Y06_lo_out[0]};
	// mantle_wire__typeBitIn16 Tile_X02_Y06_tile_id(
	// 	.in(Tile_X02_Y06_tile_id_in),
	// 	.out(Tile_X02_Y06_tile_id_out)
	// );
	// Tile_PE Tile_X02_Y07(
	// 	.SB_T0_EAST_SB_IN_B1(Tile_X03_Y07_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_IN_B16(Tile_X03_Y07_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X02_Y07_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X02_Y07_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X02_Y06_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X02_Y06_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y07_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y07_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y08_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y08_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y07_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y07_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(Tile_X01_Y07_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_IN_B16(Tile_X01_Y07_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X02_Y07_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X02_Y07_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(Tile_X03_Y07_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_IN_B16(Tile_X03_Y07_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X02_Y07_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X02_Y07_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X02_Y06_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X02_Y06_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y07_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y07_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y08_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y08_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y07_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y07_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(Tile_X01_Y07_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_IN_B16(Tile_X01_Y07_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X02_Y07_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X02_Y07_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(Tile_X03_Y07_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_IN_B16(Tile_X03_Y07_SB_T2_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X02_Y07_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X02_Y07_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X02_Y06_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X02_Y06_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y07_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y07_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y08_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y08_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y07_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y07_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(Tile_X01_Y07_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_IN_B16(Tile_X01_Y07_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X02_Y07_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X02_Y07_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X02_Y06_clk_out),
	// 	.clk_out(Tile_X02_Y07_clk_out),
	// 	.clk_pass_through(Tile_X02_Y06_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X02_Y07_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X02_Y06_config_out_config_addr),
	// 	.config_config_data(Tile_X02_Y06_config_out_config_data),
	// 	.config_out_config_addr(Tile_X02_Y07_config_out_config_addr),
	// 	.config_out_config_data(Tile_X02_Y07_config_out_config_data),
	// 	.config_out_read(Tile_X02_Y07_config_out_read),
	// 	.config_out_write(Tile_X02_Y07_config_out_write),
	// 	.config_read(Tile_X02_Y06_config_out_read),
	// 	.config_write(Tile_X02_Y06_config_out_write),
	// 	.hi(Tile_X02_Y07_hi_unq1),
	// 	.lo(Tile_X02_Y07_lo_unq1),
	// 	.read_config_data(Tile_X02_Y07_read_config_data),
	// 	.read_config_data_in(Tile_X02_Y06_read_config_data),
	// 	.reset(Tile_X02_Y06_reset_out),
	// 	.reset_out(Tile_X02_Y07_reset_out),
	// 	.stall(Tile_X02_Y06_stall_out),
	// 	.stall_out(Tile_X02_Y07_stall_out),
	// 	.tile_id(Tile_X02_Y07_tile_id_in)
	// );
	// mantle_wire__typeBit9 Tile_X02_Y07_hi(
	// 	.in(Tile_X02_Y07_hi_unq1),
	// 	.out(Tile_X02_Y07_hi_out)
	// );
	// mantle_wire__typeBit8 Tile_X02_Y07_lo(
	// 	.in(Tile_X02_Y07_lo_unq1),
	// 	.out(Tile_X02_Y07_lo_out)
	// );
	// wire [15:0] Tile_X02_Y07_tile_id_out;
	// assign Tile_X02_Y07_tile_id_out = {Tile_X02_Y07_lo_out[7], Tile_X02_Y07_lo_out[7:6], Tile_X02_Y07_lo_out[6:5], Tile_X02_Y07_lo_out[5], Tile_X02_Y07_hi_out[5], Tile_X02_Y07_lo_out[4:3], Tile_X02_Y07_lo_out[3:2], Tile_X02_Y07_lo_out[2:1], Tile_X02_Y07_hi_out[1], Tile_X02_Y07_hi_out[1:0]};
	// mantle_wire__typeBitIn16 Tile_X02_Y07_tile_id(
	// 	.in(Tile_X02_Y07_tile_id_in),
	// 	.out(Tile_X02_Y07_tile_id_out)
	// );
	// Tile_PE Tile_X02_Y08(
	// 	.SB_T0_EAST_SB_IN_B1(Tile_X03_Y08_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_IN_B16(Tile_X03_Y08_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X02_Y08_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X02_Y08_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X02_Y07_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X02_Y07_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y08_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y08_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
	// 	.SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y08_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y08_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(Tile_X01_Y08_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_IN_B16(Tile_X01_Y08_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X02_Y08_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X02_Y08_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(Tile_X03_Y08_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_IN_B16(Tile_X03_Y08_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X02_Y08_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X02_Y08_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X02_Y07_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X02_Y07_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y08_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y08_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
	// 	.SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y08_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y08_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(Tile_X01_Y08_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_IN_B16(Tile_X01_Y08_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X02_Y08_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X02_Y08_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(Tile_X03_Y08_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_IN_B16(Tile_X03_Y08_SB_T2_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X02_Y08_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X02_Y08_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X02_Y07_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X02_Y07_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y08_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y08_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
	// 	.SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y08_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y08_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(Tile_X01_Y08_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_IN_B16(Tile_X01_Y08_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X02_Y08_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X02_Y08_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X02_Y07_clk_out),
	// 	.clk_out(Tile_X02_Y08_clk_out),
	// 	.clk_pass_through(Tile_X02_Y07_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X02_Y08_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X02_Y07_config_out_config_addr),
	// 	.config_config_data(Tile_X02_Y07_config_out_config_data),
	// 	.config_out_config_addr(Tile_X02_Y08_config_out_config_addr),
	// 	.config_out_config_data(Tile_X02_Y08_config_out_config_data),
	// 	.config_out_read(Tile_X02_Y08_config_out_read),
	// 	.config_out_write(Tile_X02_Y08_config_out_write),
	// 	.config_read(Tile_X02_Y07_config_out_read),
	// 	.config_write(Tile_X02_Y07_config_out_write),
	// 	.hi(Tile_X02_Y08_hi),
	// 	.lo(Tile_X02_Y08_lo_unq1),
	// 	.read_config_data(Tile_X02_Y08_read_config_data),
	// 	.read_config_data_in(Tile_X02_Y07_read_config_data),
	// 	.reset(Tile_X02_Y07_reset_out),
	// 	.reset_out(Tile_X02_Y08_reset_out),
	// 	.stall(Tile_X02_Y07_stall_out),
	// 	.stall_out(Tile_X02_Y08_stall_out),
	// 	.tile_id(Tile_X02_Y08_tile_id_in)
	// );
	// mantle_wire__typeBit8 Tile_X02_Y08_lo(
	// 	.in(Tile_X02_Y08_lo_unq1),
	// 	.out(Tile_X02_Y08_lo_out)
	// );
	// wire [15:0] Tile_X02_Y08_tile_id_out;
	// assign Tile_X02_Y08_tile_id_out = {Tile_X02_Y08_lo_out[7], Tile_X02_Y08_lo_out[7:6], Tile_X02_Y08_lo_out[6:5], Tile_X02_Y08_lo_out[5], Tile_X02_Y08_hi[5], Tile_X02_Y08_lo_out[4:3], Tile_X02_Y08_lo_out[3:2], Tile_X02_Y08_lo_out[2], Tile_X02_Y08_hi[2], Tile_X02_Y08_lo_out[1:0], Tile_X02_Y08_lo_out[0]};
	// mantle_wire__typeBitIn16 Tile_X02_Y08_tile_id(
	// 	.in(Tile_X02_Y08_tile_id_in),
	// 	.out(Tile_X02_Y08_tile_id_out)
	// );
	// wire [15:0] Tile_X03_Y00_tile_id;
	// assign Tile_X03_Y00_tile_id = {Tile_X03_Y00_lo[7], Tile_X03_Y00_lo[7:6], Tile_X03_Y00_lo[6:5], Tile_X03_Y00_lo[5], Tile_X03_Y00_hi[5:4], Tile_X03_Y00_lo[3], Tile_X03_Y00_lo[3:2], Tile_X03_Y00_lo[2:1], Tile_X03_Y00_lo[1:0], Tile_X03_Y00_lo[0]};
	// Tile_io_core Tile_X03_Y00(
	// 	.tile_id(Tile_X03_Y00_tile_id),
	// 	.glb2io_1(glb2io_1_X03_Y00),
	// 	.f2io_1(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B1),
	// 	.io2glb_1(Tile_X03_Y00_io2glb_1),
	// 	.io2f_1(Tile_X03_Y00_io2f_1),
	// 	.glb2io_16(glb2io_16_X03_Y00),
	// 	.f2io_16(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B16),
	// 	.io2glb_16(Tile_X03_Y00_io2glb_16),
	// 	.io2f_16(Tile_X03_Y00_io2f_16),
	// 	.hi(Tile_X03_Y00_hi),
	// 	.lo(Tile_X03_Y00_lo)
	// );
	// Tile_MemCore Tile_X03_Y01(
	// 	.SB_T0_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T0_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X03_Y01_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X03_Y00_io2f_16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B16),
	// 	// .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B1),
	// 	// .SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_IN_B16(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T1_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X03_Y01_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X03_Y00_io2f_16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B16),
	// 	// .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B1),
	// 	// .SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_IN_B16(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T2_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X03_Y01_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X03_Y00_io2f_16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B16),
	// 	// .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B1),
	// 	// .SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_IN_B16(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(clk),
	// 	.clk_out(Tile_X03_Y01_clk_out),
	// 	.clk_pass_through(clk),
	// 	.clk_pass_through_out_bot(Tile_X03_Y01_clk_pass_through_out_bot),
	// 	.config_config_addr(config_3_config_addr),
	// 	.config_config_data(config_3_config_data),
	// 	.config_out_config_addr(Tile_X03_Y01_config_out_config_addr),
	// 	.config_out_config_data(Tile_X03_Y01_config_out_config_data),
	// 	.config_out_read(Tile_X03_Y01_config_out_read),
	// 	.config_out_write(Tile_X03_Y01_config_out_write),
	// 	.config_read(config_3_read),
	// 	.config_write(config_3_write),
	// 	.hi(Tile_X03_Y01_hi_unq1),
	// 	.lo(Tile_X03_Y01_lo_unq1),
	// 	.read_config_data(Tile_X03_Y01_read_config_data),
	// 	.read_config_data_in(const_0_32_out),
	// 	.reset(reset),
	// 	.reset_out(Tile_X03_Y01_reset_out),
	// 	.stall(stall[3]),
	// 	.stall_out(Tile_X03_Y01_stall_out),
	// 	.tile_id(Tile_X03_Y01_tile_id_in)
	// );
	// mantle_wire__typeBit9 Tile_X03_Y01_hi(
	// 	.in(Tile_X03_Y01_hi_unq1),
	// 	.out(Tile_X03_Y01_hi_out)
	// );
	// mantle_wire__typeBit8 Tile_X03_Y01_lo(
	// 	.in(Tile_X03_Y01_lo_unq1),
	// 	.out(Tile_X03_Y01_lo_out)
	// );
	// wire [15:0] Tile_X03_Y01_tile_id_out;
	// assign Tile_X03_Y01_tile_id_out = {Tile_X03_Y01_lo_out[7], Tile_X03_Y01_lo_out[7:6], Tile_X03_Y01_lo_out[6:5], Tile_X03_Y01_lo_out[5], Tile_X03_Y01_hi_out[5:4], Tile_X03_Y01_lo_out[3], Tile_X03_Y01_lo_out[3:2], Tile_X03_Y01_lo_out[2:1], Tile_X03_Y01_lo_out[1:0], Tile_X03_Y01_hi_out[0]};
	// mantle_wire__typeBitIn16 Tile_X03_Y01_tile_id(
	// 	.in(Tile_X03_Y01_tile_id_in),
	// 	.out(Tile_X03_Y01_tile_id_out)
	// );
	// Tile_PE Tile_X03_Y02(
	// 	.SB_T0_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T0_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X03_Y02_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B16),
	// 	// .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B1),
	// 	// .SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B16),
	// 	// .SB_T0_WEST_SB_IN_B1(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B1),
	// 	// .SB_T0_WEST_SB_IN_B16(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T1_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X03_Y02_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B16),
	// 	// .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B1),
	// 	// .SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B16),
	// 	// .SB_T1_WEST_SB_IN_B1(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B1),
	// 	// .SB_T1_WEST_SB_IN_B16(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T2_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X03_Y02_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B16),
	// 	// .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B1),
	// 	// .SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B16),
	// 	// .SB_T2_WEST_SB_IN_B1(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B1),
	// 	// .SB_T2_WEST_SB_IN_B16(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X03_Y01_clk_out),
	// 	.clk_out(Tile_X03_Y02_clk_out),
	// 	.clk_pass_through(Tile_X03_Y01_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X03_Y02_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X03_Y01_config_out_config_addr),
	// 	.config_config_data(Tile_X03_Y01_config_out_config_data),
	// 	.config_out_config_addr(Tile_X03_Y02_config_out_config_addr),
	// 	.config_out_config_data(Tile_X03_Y02_config_out_config_data),
	// 	.config_out_read(Tile_X03_Y02_config_out_read),
	// 	.config_out_write(Tile_X03_Y02_config_out_write),
	// 	.config_read(Tile_X03_Y01_config_out_read),
	// 	.config_write(Tile_X03_Y01_config_out_write),
	// 	.hi(Tile_X03_Y02_hi_unq1),
	// 	.lo(Tile_X03_Y02_lo_unq1),
	// 	.read_config_data(Tile_X03_Y02_read_config_data),
	// 	.read_config_data_in(Tile_X03_Y01_read_config_data),
	// 	.reset(Tile_X03_Y01_reset_out),
	// 	.reset_out(Tile_X03_Y02_reset_out),
	// 	.stall(Tile_X03_Y01_stall_out),
	// 	.stall_out(Tile_X03_Y02_stall_out),
	// 	.tile_id(Tile_X03_Y02_tile_id_in)
	// );
	// mantle_wire__typeBit9 Tile_X03_Y02_hi(
	// 	.in(Tile_X03_Y02_hi_unq1),
	// 	.out(Tile_X03_Y02_hi_out)
	// );
	// mantle_wire__typeBit8 Tile_X03_Y02_lo(
	// 	.in(Tile_X03_Y02_lo_unq1),
	// 	.out(Tile_X03_Y02_lo_out)
	// );
	// wire [15:0] Tile_X03_Y02_tile_id_out;
	// assign Tile_X03_Y02_tile_id_out = {Tile_X03_Y02_lo_out[7], Tile_X03_Y02_lo_out[7:6], Tile_X03_Y02_lo_out[6:5], Tile_X03_Y02_lo_out[5], Tile_X03_Y02_hi_out[5:4], Tile_X03_Y02_lo_out[3], Tile_X03_Y02_lo_out[3:2], Tile_X03_Y02_lo_out[2:1], Tile_X03_Y02_lo_out[1], Tile_X03_Y02_hi_out[1], Tile_X03_Y02_lo_out[0]};
	// mantle_wire__typeBitIn16 Tile_X03_Y02_tile_id(
	// 	.in(Tile_X03_Y02_tile_id_in),
	// 	.out(Tile_X03_Y02_tile_id_out)
	// );
	// Tile_PE Tile_X03_Y03(
	// 	.SB_T0_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T0_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X03_Y03_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_IN_B16(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T1_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X03_Y03_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_IN_B16(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T2_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X03_Y03_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_IN_B16(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X03_Y02_clk_out),
	// 	.clk_out(Tile_X03_Y03_clk_out),
	// 	.clk_pass_through(Tile_X03_Y02_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X03_Y03_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X03_Y02_config_out_config_addr),
	// 	.config_config_data(Tile_X03_Y02_config_out_config_data),
	// 	.config_out_config_addr(Tile_X03_Y03_config_out_config_addr),
	// 	.config_out_config_data(Tile_X03_Y03_config_out_config_data),
	// 	.config_out_read(Tile_X03_Y03_config_out_read),
	// 	.config_out_write(Tile_X03_Y03_config_out_write),
	// 	.config_read(Tile_X03_Y02_config_out_read),
	// 	.config_write(Tile_X03_Y02_config_out_write),
	// 	.hi(Tile_X03_Y03_hi_unq1),
	// 	.lo(Tile_X03_Y03_lo_unq1),
	// 	.read_config_data(Tile_X03_Y03_read_config_data),
	// 	.read_config_data_in(Tile_X03_Y02_read_config_data),
	// 	.reset(Tile_X03_Y02_reset_out),
	// 	.reset_out(Tile_X03_Y03_reset_out),
	// 	.stall(Tile_X03_Y02_stall_out),
	// 	.stall_out(Tile_X03_Y03_stall_out),
	// 	.tile_id(Tile_X03_Y03_tile_id_in)
	// );
	// mantle_wire__typeBit9 Tile_X03_Y03_hi(
	// 	.in(Tile_X03_Y03_hi_unq1),
	// 	.out(Tile_X03_Y03_hi_out)
	// );
	// mantle_wire__typeBit8 Tile_X03_Y03_lo(
	// 	.in(Tile_X03_Y03_lo_unq1),
	// 	.out(Tile_X03_Y03_lo_out)
	// );
	// wire [15:0] Tile_X03_Y03_tile_id_out;
	// assign Tile_X03_Y03_tile_id_out = {Tile_X03_Y03_lo_out[7], Tile_X03_Y03_lo_out[7:6], Tile_X03_Y03_lo_out[6:5], Tile_X03_Y03_lo_out[5], Tile_X03_Y03_hi_out[5:4], Tile_X03_Y03_lo_out[3], Tile_X03_Y03_lo_out[3:2], Tile_X03_Y03_lo_out[2:1], Tile_X03_Y03_lo_out[1], Tile_X03_Y03_hi_out[1:0]};
	// mantle_wire__typeBitIn16 Tile_X03_Y03_tile_id(
	// 	.in(Tile_X03_Y03_tile_id_in),
	// 	.out(Tile_X03_Y03_tile_id_out)
	// );
	// Tile_PE Tile_X03_Y04(
	// 	.SB_T0_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T0_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X03_Y04_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y05_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y05_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_IN_B16(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T1_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X03_Y04_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y05_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y05_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_IN_B16(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T2_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X03_Y04_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y05_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y05_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_IN_B16(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X03_Y03_clk_out),
	// 	.clk_out(Tile_X03_Y04_clk_out),
	// 	.clk_pass_through(Tile_X03_Y03_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X03_Y04_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X03_Y03_config_out_config_addr),
	// 	.config_config_data(Tile_X03_Y03_config_out_config_data),
	// 	.config_out_config_addr(Tile_X03_Y04_config_out_config_addr),
	// 	.config_out_config_data(Tile_X03_Y04_config_out_config_data),
	// 	.config_out_read(Tile_X03_Y04_config_out_read),
	// 	.config_out_write(Tile_X03_Y04_config_out_write),
	// 	.config_read(Tile_X03_Y03_config_out_read),
	// 	.config_write(Tile_X03_Y03_config_out_write),
	// 	.hi(Tile_X03_Y04_hi_unq1),
	// 	.lo(Tile_X03_Y04_lo_unq1),
	// 	.read_config_data(Tile_X03_Y04_read_config_data),
	// 	.read_config_data_in(Tile_X03_Y03_read_config_data),
	// 	.reset(Tile_X03_Y03_reset_out),
	// 	.reset_out(Tile_X03_Y04_reset_out),
	// 	.stall(Tile_X03_Y03_stall_out),
	// 	.stall_out(Tile_X03_Y04_stall_out),
	// 	.tile_id(Tile_X03_Y04_tile_id_in)
	// );
	// mantle_wire__typeBit9 Tile_X03_Y04_hi(
	// 	.in(Tile_X03_Y04_hi_unq1),
	// 	.out(Tile_X03_Y04_hi_out)
	// );
	// mantle_wire__typeBit8 Tile_X03_Y04_lo(
	// 	.in(Tile_X03_Y04_lo_unq1),
	// 	.out(Tile_X03_Y04_lo_out)
	// );
	// wire [15:0] Tile_X03_Y04_tile_id_out;
	// assign Tile_X03_Y04_tile_id_out = {Tile_X03_Y04_lo_out[7], Tile_X03_Y04_lo_out[7:6], Tile_X03_Y04_lo_out[6:5], Tile_X03_Y04_lo_out[5], Tile_X03_Y04_hi_out[5:4], Tile_X03_Y04_lo_out[3], Tile_X03_Y04_lo_out[3:2], Tile_X03_Y04_lo_out[2:1], Tile_X03_Y04_hi_out[1], Tile_X03_Y04_lo_out[0], Tile_X03_Y04_lo_out[0]};
	// mantle_wire__typeBitIn16 Tile_X03_Y04_tile_id(
	// 	.in(Tile_X03_Y04_tile_id_in),
	// 	.out(Tile_X03_Y04_tile_id_out)
	// );
	// Tile_MemCore Tile_X03_Y05(
	// 	.SB_T0_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T0_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X03_Y05_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X03_Y05_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y05_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y05_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y06_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y06_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y05_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y05_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(Tile_X02_Y05_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_IN_B16(Tile_X02_Y05_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X03_Y05_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X03_Y05_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T1_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X03_Y05_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X03_Y05_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y05_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y05_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y06_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y06_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y05_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y05_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(Tile_X02_Y05_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_IN_B16(Tile_X02_Y05_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X03_Y05_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X03_Y05_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T2_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X03_Y05_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X03_Y05_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y05_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y05_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y06_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y06_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y05_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y05_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(Tile_X02_Y05_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_IN_B16(Tile_X02_Y05_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X03_Y05_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X03_Y05_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X03_Y04_clk_out),
	// 	.clk_out(Tile_X03_Y05_clk_out),
	// 	.clk_pass_through(Tile_X03_Y04_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X03_Y05_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X03_Y04_config_out_config_addr),
	// 	.config_config_data(Tile_X03_Y04_config_out_config_data),
	// 	.config_out_config_addr(Tile_X03_Y05_config_out_config_addr),
	// 	.config_out_config_data(Tile_X03_Y05_config_out_config_data),
	// 	.config_out_read(Tile_X03_Y05_config_out_read),
	// 	.config_out_write(Tile_X03_Y05_config_out_write),
	// 	.config_read(Tile_X03_Y04_config_out_read),
	// 	.config_write(Tile_X03_Y04_config_out_write),
	// 	.hi(Tile_X03_Y05_hi_unq1),
	// 	.lo(Tile_X03_Y05_lo_unq1),
	// 	.read_config_data(Tile_X03_Y05_read_config_data),
	// 	.read_config_data_in(Tile_X03_Y04_read_config_data),
	// 	.reset(Tile_X03_Y04_reset_out),
	// 	.reset_out(Tile_X03_Y05_reset_out),
	// 	.stall(Tile_X03_Y04_stall_out),
	// 	.stall_out(Tile_X03_Y05_stall_out),
	// 	.tile_id(Tile_X03_Y05_tile_id_in)
	// );
	// mantle_wire__typeBit9 Tile_X03_Y05_hi(
	// 	.in(Tile_X03_Y05_hi_unq1),
	// 	.out(Tile_X03_Y05_hi_out)
	// );
	// mantle_wire__typeBit8 Tile_X03_Y05_lo(
	// 	.in(Tile_X03_Y05_lo_unq1),
	// 	.out(Tile_X03_Y05_lo_out)
	// );
	// wire [15:0] Tile_X03_Y05_tile_id_out;
	// assign Tile_X03_Y05_tile_id_out = {Tile_X03_Y05_lo_out[7], Tile_X03_Y05_lo_out[7:6], Tile_X03_Y05_lo_out[6:5], Tile_X03_Y05_lo_out[5], Tile_X03_Y05_hi_out[5:4], Tile_X03_Y05_lo_out[3], Tile_X03_Y05_lo_out[3:2], Tile_X03_Y05_lo_out[2:1], Tile_X03_Y05_hi_out[1], Tile_X03_Y05_lo_out[0], Tile_X03_Y05_hi_out[0]};
	// mantle_wire__typeBitIn16 Tile_X03_Y05_tile_id(
	// 	.in(Tile_X03_Y05_tile_id_in),
	// 	.out(Tile_X03_Y05_tile_id_out)
	// );
	// Tile_PE Tile_X03_Y06(
	// 	.SB_T0_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T0_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X03_Y06_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X03_Y06_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X03_Y05_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X03_Y05_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y06_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y06_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y07_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y07_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y06_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y06_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(Tile_X02_Y06_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_IN_B16(Tile_X02_Y06_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X03_Y06_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X03_Y06_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T1_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X03_Y06_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X03_Y06_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X03_Y05_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X03_Y05_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y06_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y06_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y07_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y07_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y06_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y06_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(Tile_X02_Y06_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_IN_B16(Tile_X02_Y06_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X03_Y06_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X03_Y06_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T2_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X03_Y06_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X03_Y06_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X03_Y05_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X03_Y05_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y06_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y06_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y07_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y07_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y06_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y06_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(Tile_X02_Y06_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_IN_B16(Tile_X02_Y06_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X03_Y06_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X03_Y06_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X03_Y05_clk_out),
	// 	.clk_out(Tile_X03_Y06_clk_out),
	// 	.clk_pass_through(Tile_X03_Y05_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X03_Y06_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X03_Y05_config_out_config_addr),
	// 	.config_config_data(Tile_X03_Y05_config_out_config_data),
	// 	.config_out_config_addr(Tile_X03_Y06_config_out_config_addr),
	// 	.config_out_config_data(Tile_X03_Y06_config_out_config_data),
	// 	.config_out_read(Tile_X03_Y06_config_out_read),
	// 	.config_out_write(Tile_X03_Y06_config_out_write),
	// 	.config_read(Tile_X03_Y05_config_out_read),
	// 	.config_write(Tile_X03_Y05_config_out_write),
	// 	.hi(Tile_X03_Y06_hi_unq1),
	// 	.lo(Tile_X03_Y06_lo_unq1),
	// 	.read_config_data(Tile_X03_Y06_read_config_data),
	// 	.read_config_data_in(Tile_X03_Y05_read_config_data),
	// 	.reset(Tile_X03_Y05_reset_out),
	// 	.reset_out(Tile_X03_Y06_reset_out),
	// 	.stall(Tile_X03_Y05_stall_out),
	// 	.stall_out(Tile_X03_Y06_stall_out),
	// 	.tile_id(Tile_X03_Y06_tile_id_in)
	// );
	// mantle_wire__typeBit9 Tile_X03_Y06_hi(
	// 	.in(Tile_X03_Y06_hi_unq1),
	// 	.out(Tile_X03_Y06_hi_out)
	// );
	// mantle_wire__typeBit8 Tile_X03_Y06_lo(
	// 	.in(Tile_X03_Y06_lo_unq1),
	// 	.out(Tile_X03_Y06_lo_out)
	// );
	// wire [15:0] Tile_X03_Y06_tile_id_out;
	// assign Tile_X03_Y06_tile_id_out = {Tile_X03_Y06_lo_out[7], Tile_X03_Y06_lo_out[7:6], Tile_X03_Y06_lo_out[6:5], Tile_X03_Y06_lo_out[5], Tile_X03_Y06_hi_out[5:4], Tile_X03_Y06_lo_out[3], Tile_X03_Y06_lo_out[3:2], Tile_X03_Y06_lo_out[2:1], Tile_X03_Y06_hi_out[1], Tile_X03_Y06_hi_out[1], Tile_X03_Y06_lo_out[0]};
	// mantle_wire__typeBitIn16 Tile_X03_Y06_tile_id(
	// 	.in(Tile_X03_Y06_tile_id_in),
	// 	.out(Tile_X03_Y06_tile_id_out)
	// );
	// Tile_PE Tile_X03_Y07(
	// 	.SB_T0_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T0_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X03_Y07_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X03_Y07_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X03_Y06_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X03_Y06_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y07_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y07_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y08_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y08_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y07_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y07_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(Tile_X02_Y07_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_IN_B16(Tile_X02_Y07_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X03_Y07_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X03_Y07_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T1_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X03_Y07_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X03_Y07_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X03_Y06_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X03_Y06_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y07_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y07_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y08_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y08_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y07_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y07_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(Tile_X02_Y07_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_IN_B16(Tile_X02_Y07_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X03_Y07_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X03_Y07_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T2_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X03_Y07_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X03_Y07_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X03_Y06_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X03_Y06_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y07_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y07_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y08_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y08_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y07_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y07_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(Tile_X02_Y07_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_IN_B16(Tile_X02_Y07_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X03_Y07_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X03_Y07_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X03_Y06_clk_out),
	// 	.clk_out(Tile_X03_Y07_clk_out),
	// 	.clk_pass_through(Tile_X03_Y06_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X03_Y07_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X03_Y06_config_out_config_addr),
	// 	.config_config_data(Tile_X03_Y06_config_out_config_data),
	// 	.config_out_config_addr(Tile_X03_Y07_config_out_config_addr),
	// 	.config_out_config_data(Tile_X03_Y07_config_out_config_data),
	// 	.config_out_read(Tile_X03_Y07_config_out_read),
	// 	.config_out_write(Tile_X03_Y07_config_out_write),
	// 	.config_read(Tile_X03_Y06_config_out_read),
	// 	.config_write(Tile_X03_Y06_config_out_write),
	// 	.hi(Tile_X03_Y07_hi_unq1),
	// 	.lo(Tile_X03_Y07_lo_unq1),
	// 	.read_config_data(Tile_X03_Y07_read_config_data),
	// 	.read_config_data_in(Tile_X03_Y06_read_config_data),
	// 	.reset(Tile_X03_Y06_reset_out),
	// 	.reset_out(Tile_X03_Y07_reset_out),
	// 	.stall(Tile_X03_Y06_stall_out),
	// 	.stall_out(Tile_X03_Y07_stall_out),
	// 	.tile_id(Tile_X03_Y07_tile_id_in)
	// );
	// mantle_wire__typeBit9 Tile_X03_Y07_hi(
	// 	.in(Tile_X03_Y07_hi_unq1),
	// 	.out(Tile_X03_Y07_hi_out)
	// );
	// mantle_wire__typeBit8 Tile_X03_Y07_lo(
	// 	.in(Tile_X03_Y07_lo_unq1),
	// 	.out(Tile_X03_Y07_lo_out)
	// );
	// wire [15:0] Tile_X03_Y07_tile_id_out;
	// assign Tile_X03_Y07_tile_id_out = {Tile_X03_Y07_lo_out[7], Tile_X03_Y07_lo_out[7:6], Tile_X03_Y07_lo_out[6:5], Tile_X03_Y07_lo_out[5], Tile_X03_Y07_hi_out[5:4], Tile_X03_Y07_lo_out[3], Tile_X03_Y07_lo_out[3:2], Tile_X03_Y07_lo_out[2:1], Tile_X03_Y07_hi_out[1], Tile_X03_Y07_hi_out[1:0]};
	// mantle_wire__typeBitIn16 Tile_X03_Y07_tile_id(
	// 	.in(Tile_X03_Y07_tile_id_in),
	// 	.out(Tile_X03_Y07_tile_id_out)
	// );
	// Tile_PE Tile_X03_Y08(
	// 	.SB_T0_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T0_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T0_EAST_SB_OUT_B1(Tile_X03_Y08_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_EAST_SB_OUT_B16(Tile_X03_Y08_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_IN_B1(Tile_X03_Y07_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_IN_B16(Tile_X03_Y07_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y08_SB_T0_NORTH_SB_OUT_B1),
	// 	.SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y08_SB_T0_NORTH_SB_OUT_B16),
	// 	.SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
	// 	.SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
	// 	.SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y08_SB_T0_SOUTH_SB_OUT_B1),
	// 	.SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y08_SB_T0_SOUTH_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_IN_B1(Tile_X02_Y08_SB_T0_EAST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_IN_B16(Tile_X02_Y08_SB_T0_EAST_SB_OUT_B16),
	// 	.SB_T0_WEST_SB_OUT_B1(Tile_X03_Y08_SB_T0_WEST_SB_OUT_B1),
	// 	.SB_T0_WEST_SB_OUT_B16(Tile_X03_Y08_SB_T0_WEST_SB_OUT_B16),
	// 	.SB_T1_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T1_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T1_EAST_SB_OUT_B1(Tile_X03_Y08_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_EAST_SB_OUT_B16(Tile_X03_Y08_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_IN_B1(Tile_X03_Y07_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_IN_B16(Tile_X03_Y07_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y08_SB_T1_NORTH_SB_OUT_B1),
	// 	.SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y08_SB_T1_NORTH_SB_OUT_B16),
	// 	.SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
	// 	.SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
	// 	.SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y08_SB_T1_SOUTH_SB_OUT_B1),
	// 	.SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y08_SB_T1_SOUTH_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_IN_B1(Tile_X02_Y08_SB_T1_EAST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_IN_B16(Tile_X02_Y08_SB_T1_EAST_SB_OUT_B16),
	// 	.SB_T1_WEST_SB_OUT_B1(Tile_X03_Y08_SB_T1_WEST_SB_OUT_B1),
	// 	.SB_T1_WEST_SB_OUT_B16(Tile_X03_Y08_SB_T1_WEST_SB_OUT_B16),
	// 	.SB_T2_EAST_SB_IN_B1(const_0_1_out),
	// 	.SB_T2_EAST_SB_IN_B16(const_0_16_out),
	// 	.SB_T2_EAST_SB_OUT_B1(Tile_X03_Y08_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_EAST_SB_OUT_B16(Tile_X03_Y08_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_IN_B1(Tile_X03_Y07_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_IN_B16(Tile_X03_Y07_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y08_SB_T2_NORTH_SB_OUT_B1),
	// 	.SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y08_SB_T2_NORTH_SB_OUT_B16),
	// 	.SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
	// 	.SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
	// 	.SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y08_SB_T2_SOUTH_SB_OUT_B1),
	// 	.SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y08_SB_T2_SOUTH_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_IN_B1(Tile_X02_Y08_SB_T2_EAST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_IN_B16(Tile_X02_Y08_SB_T2_EAST_SB_OUT_B16),
	// 	.SB_T2_WEST_SB_OUT_B1(Tile_X03_Y08_SB_T2_WEST_SB_OUT_B1),
	// 	.SB_T2_WEST_SB_OUT_B16(Tile_X03_Y08_SB_T2_WEST_SB_OUT_B16),
	// 	.clk(Tile_X03_Y07_clk_out),
	// 	.clk_out(Tile_X03_Y08_clk_out),
	// 	.clk_pass_through(Tile_X03_Y07_clk_pass_through_out_bot),
	// 	.clk_pass_through_out_bot(Tile_X03_Y08_clk_pass_through_out_bot),
	// 	.config_config_addr(Tile_X03_Y07_config_out_config_addr),
	// 	.config_config_data(Tile_X03_Y07_config_out_config_data),
	// 	.config_out_config_addr(Tile_X03_Y08_config_out_config_addr),
	// 	.config_out_config_data(Tile_X03_Y08_config_out_config_data),
	// 	.config_out_read(Tile_X03_Y08_config_out_read),
	// 	.config_out_write(Tile_X03_Y08_config_out_write),
	// 	.config_read(Tile_X03_Y07_config_out_read),
	// 	.config_write(Tile_X03_Y07_config_out_write),
	// 	.hi(Tile_X03_Y08_hi_unq1),
	// 	.lo(Tile_X03_Y08_lo_unq1),
	// 	.read_config_data(Tile_X03_Y08_read_config_data),
	// 	.read_config_data_in(Tile_X03_Y07_read_config_data),
	// 	.reset(Tile_X03_Y07_reset_out),
	// 	.reset_out(Tile_X03_Y08_reset_out),
	// 	.stall(Tile_X03_Y07_stall_out),
	// 	.stall_out(Tile_X03_Y08_stall_out),
	// 	.tile_id(Tile_X03_Y08_tile_id_in)
	// );
	// mantle_wire__typeBit9 Tile_X03_Y08_hi(
	// 	.in(Tile_X03_Y08_hi_unq1),
	// 	.out(Tile_X03_Y08_hi_out)
	// );
	// mantle_wire__typeBit8 Tile_X03_Y08_lo(
	// 	.in(Tile_X03_Y08_lo_unq1),
	// 	.out(Tile_X03_Y08_lo_out)
	// );
	// wire [15:0] Tile_X03_Y08_tile_id_out;
	// assign Tile_X03_Y08_tile_id_out = {Tile_X03_Y08_lo_out[7], Tile_X03_Y08_lo_out[7:6], Tile_X03_Y08_lo_out[6:5], Tile_X03_Y08_lo_out[5], Tile_X03_Y08_hi_out[5:4], Tile_X03_Y08_lo_out[3], Tile_X03_Y08_lo_out[3:2], Tile_X03_Y08_lo_out[2], Tile_X03_Y08_hi_out[2], Tile_X03_Y08_lo_out[1:0], Tile_X03_Y08_lo_out[0]};
	// mantle_wire__typeBitIn16 Tile_X03_Y08_tile_id(
	// 	.in(Tile_X03_Y08_tile_id_in),
	// 	.out(Tile_X03_Y08_tile_id_out)
	// );
	coreir_const #(
		.value(1'h0),
		.width(1)
	) const_0_1(.out(const_0_1_out));
	coreir_const #(
		.value(16'h0000),
		.width(16)
	) const_0_16(.out(const_0_16_out));
	coreir_const #(
		.value(32'h00000000),
		.width(32)
	) const_0_32(.out(const_0_32_out));

	// Change to the End line (Current should change to Y02)
	Or4x32 read_config_data_or_final(
		.I0(Tile_X00_Y02_read_config_data),	// Only connected with One PE for Tile_X00_Y02
		.I1(Tile_X01_Y02_read_config_data),
		// .I2(Tile_X02_Y02_read_config_data),
		// .I3(Tile_X03_Y02_read_config_data),
		.O(read_config_data_or_final_O)
	);
	assign io2glb_16_X00_Y00 = Tile_X00_Y00_io2glb_16;
	assign io2glb_16_X01_Y00 = Tile_X01_Y00_io2glb_16;
	// assign io2glb_16_X02_Y00 = Tile_X02_Y00_io2glb_16;
	// assign io2glb_16_X03_Y00 = Tile_X03_Y00_io2glb_16;
	assign io2glb_1_X00_Y00 = Tile_X00_Y00_io2glb_1;
	assign io2glb_1_X01_Y00 = Tile_X01_Y00_io2glb_1;
	// assign io2glb_1_X02_Y00 = Tile_X02_Y00_io2glb_1;
	// assign io2glb_1_X03_Y00 = Tile_X03_Y00_io2glb_1;
	assign read_config_data = read_config_data_or_final_O;
endmodule
module Garnet (
	clk,
	config_0_config_addr,
	config_0_config_data,
	config_0_read,
	config_0_write,
	config_1_config_addr,
	config_1_config_data,
	config_1_read,
	config_1_write,
	config_2_config_addr,
	config_2_config_data,
	config_2_read,
	config_2_write,
	config_3_config_addr,
	config_3_config_data,
	config_3_read,
	config_3_write,
	glb2io_16_X00_Y00,
	glb2io_16_X01_Y00,
	// glb2io_16_X02_Y00,
	// glb2io_16_X03_Y00,
	glb2io_1_X00_Y00,
	glb2io_1_X01_Y00,
	// glb2io_1_X02_Y00,
	// glb2io_1_X03_Y00,
	io2glb_16_X00_Y00,
	io2glb_16_X01_Y00,
	// io2glb_16_X02_Y00,
	// io2glb_16_X03_Y00,
	io2glb_1_X00_Y00,
	io2glb_1_X01_Y00,
	// io2glb_1_X02_Y00,
	// io2glb_1_X03_Y00,
	read_config_data,
	reset,
	stall
);
	input clk;
	input [31:0] config_0_config_addr;
	input [31:0] config_0_config_data;
	input [0:0] config_0_read;
	input [0:0] config_0_write;
	input [31:0] config_1_config_addr;
	input [31:0] config_1_config_data;
	input [0:0] config_1_read;
	input [0:0] config_1_write;
	input [31:0] config_2_config_addr;
	input [31:0] config_2_config_data;
	input [0:0] config_2_read;
	input [0:0] config_2_write;
	input [31:0] config_3_config_addr;
	input [31:0] config_3_config_data;
	input [0:0] config_3_read;
	input [0:0] config_3_write;
	input [15:0] glb2io_16_X00_Y00;
	input [15:0] glb2io_16_X01_Y00;
	// input [15:0] glb2io_16_X02_Y00;
	// input [15:0] glb2io_16_X03_Y00;
	input [0:0] glb2io_1_X00_Y00;
	input [0:0] glb2io_1_X01_Y00;
	// input [0:0] glb2io_1_X02_Y00;
	// input [0:0] glb2io_1_X03_Y00;
	output [15:0] io2glb_16_X00_Y00;
	output [15:0] io2glb_16_X01_Y00;
	// output [15:0] io2glb_16_X02_Y00;
	// output [15:0] io2glb_16_X03_Y00;
	output [0:0] io2glb_1_X00_Y00;
	output [0:0] io2glb_1_X01_Y00;
	// output [0:0] io2glb_1_X02_Y00;
	// output [0:0] io2glb_1_X03_Y00;
	output [31:0] read_config_data;
	input reset;
	input [3:0] stall;
	wire [15:0] Interconnect_inst0_io2glb_16_X00_Y00;
	wire [15:0] Interconnect_inst0_io2glb_16_X01_Y00;
	// wire [15:0] Interconnect_inst0_io2glb_16_X02_Y00;
	// wire [15:0] Interconnect_inst0_io2glb_16_X03_Y00;
	wire [0:0] Interconnect_inst0_io2glb_1_X00_Y00;
	wire [0:0] Interconnect_inst0_io2glb_1_X01_Y00;
	// wire [0:0] Interconnect_inst0_io2glb_1_X02_Y00;
	// wire [0:0] Interconnect_inst0_io2glb_1_X03_Y00;
	wire [31:0] Interconnect_inst0_read_config_data;
	Interconnect Interconnect_inst0(
		.clk(clk),
		.config_0_config_addr(config_0_config_addr),
		.config_0_config_data(config_0_config_data),
		.config_0_read(config_0_read),
		.config_0_write(config_0_write),
		.config_1_config_addr(config_1_config_addr),
		.config_1_config_data(config_1_config_data),
		.config_1_read(config_1_read),
		.config_1_write(config_1_write),
		.config_2_config_addr(config_2_config_addr),
		.config_2_config_data(config_2_config_data),
		.config_2_read(config_2_read),
		.config_2_write(config_2_write),
		.config_3_config_addr(config_3_config_addr),
		.config_3_config_data(config_3_config_data),
		.config_3_read(config_3_read),
		.config_3_write(config_3_write),
		.glb2io_16_X00_Y00(glb2io_16_X00_Y00),
		.glb2io_16_X01_Y00(glb2io_16_X01_Y00),
		// .glb2io_16_X02_Y00(glb2io_16_X02_Y00),
		// .glb2io_16_X03_Y00(glb2io_16_X03_Y00),
		.glb2io_1_X00_Y00(glb2io_1_X00_Y00),
		.glb2io_1_X01_Y00(glb2io_1_X01_Y00),
		// .glb2io_1_X02_Y00(glb2io_1_X02_Y00),
		// .glb2io_1_X03_Y00(glb2io_1_X03_Y00),
		.io2glb_16_X00_Y00(Interconnect_inst0_io2glb_16_X00_Y00),
		.io2glb_16_X01_Y00(Interconnect_inst0_io2glb_16_X01_Y00),
		// .io2glb_16_X02_Y00(Interconnect_inst0_io2glb_16_X02_Y00),
		// .io2glb_16_X03_Y00(Interconnect_inst0_io2glb_16_X03_Y00),
		.io2glb_1_X00_Y00(Interconnect_inst0_io2glb_1_X00_Y00),
		.io2glb_1_X01_Y00(Interconnect_inst0_io2glb_1_X01_Y00),
		// .io2glb_1_X02_Y00(Interconnect_inst0_io2glb_1_X02_Y00),
		// .io2glb_1_X03_Y00(Interconnect_inst0_io2glb_1_X03_Y00),
		.read_config_data(Interconnect_inst0_read_config_data),
		.reset(reset),
		.stall(stall)
	);
	assign io2glb_16_X00_Y00 = Interconnect_inst0_io2glb_16_X00_Y00;
	assign io2glb_16_X01_Y00 = Interconnect_inst0_io2glb_16_X01_Y00;
	// assign io2glb_16_X02_Y00 = Interconnect_inst0_io2glb_16_X02_Y00;
	// assign io2glb_16_X03_Y00 = Interconnect_inst0_io2glb_16_X03_Y00;
	assign io2glb_1_X00_Y00 = Interconnect_inst0_io2glb_1_X00_Y00;
	assign io2glb_1_X01_Y00 = Interconnect_inst0_io2glb_1_X01_Y00;
	// assign io2glb_1_X02_Y00 = Interconnect_inst0_io2glb_1_X02_Y00;
	// assign io2glb_1_X03_Y00 = Interconnect_inst0_io2glb_1_X03_Y00;
	assign read_config_data = Interconnect_inst0_read_config_data;
endmodule
